magic
tech gf180mcuD
magscale 1 10
timestamp 1701795194
<< metal1 >>
rect 53778 56590 53790 56642
rect 53842 56639 53854 56642
rect 55010 56639 55022 56642
rect 53842 56593 55022 56639
rect 53842 56590 53854 56593
rect 55010 56590 55022 56593
rect 55074 56590 55086 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 10334 56306 10386 56318
rect 10334 56242 10386 56254
rect 11006 56306 11058 56318
rect 11006 56242 11058 56254
rect 13694 56306 13746 56318
rect 13694 56242 13746 56254
rect 25230 56306 25282 56318
rect 25230 56242 25282 56254
rect 34302 56306 34354 56318
rect 34302 56242 34354 56254
rect 48974 56306 49026 56318
rect 48974 56242 49026 56254
rect 52222 56306 52274 56318
rect 52222 56242 52274 56254
rect 54126 56306 54178 56318
rect 54126 56242 54178 56254
rect 55022 56306 55074 56318
rect 55022 56242 55074 56254
rect 55470 56306 55522 56318
rect 55470 56242 55522 56254
rect 33742 56194 33794 56206
rect 33742 56130 33794 56142
rect 25118 56082 25170 56094
rect 32286 56082 32338 56094
rect 31154 56030 31166 56082
rect 31218 56030 31230 56082
rect 25118 56018 25170 56030
rect 32286 56018 32338 56030
rect 33294 56082 33346 56094
rect 33294 56018 33346 56030
rect 33854 56082 33906 56094
rect 48178 56030 48190 56082
rect 48242 56030 48254 56082
rect 51202 56030 51214 56082
rect 51266 56030 51278 56082
rect 33854 56018 33906 56030
rect 8318 55970 8370 55982
rect 8318 55906 8370 55918
rect 19182 55970 19234 55982
rect 19182 55906 19234 55918
rect 25790 55970 25842 55982
rect 25790 55906 25842 55918
rect 26910 55970 26962 55982
rect 33518 55970 33570 55982
rect 55918 55970 55970 55982
rect 29586 55918 29598 55970
rect 29650 55918 29662 55970
rect 34738 55918 34750 55970
rect 34802 55918 34814 55970
rect 26910 55906 26962 55918
rect 33518 55906 33570 55918
rect 55918 55906 55970 55918
rect 25230 55858 25282 55870
rect 25230 55794 25282 55806
rect 58158 55858 58210 55870
rect 58158 55794 58210 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 48190 55522 48242 55534
rect 48190 55458 48242 55470
rect 49646 55410 49698 55422
rect 29362 55358 29374 55410
rect 29426 55358 29438 55410
rect 49646 55346 49698 55358
rect 53678 55410 53730 55422
rect 53678 55346 53730 55358
rect 33742 55298 33794 55310
rect 23762 55246 23774 55298
rect 23826 55246 23838 55298
rect 29698 55246 29710 55298
rect 29762 55246 29774 55298
rect 33058 55246 33070 55298
rect 33122 55246 33134 55298
rect 33742 55234 33794 55246
rect 34078 55298 34130 55310
rect 36990 55298 37042 55310
rect 39566 55298 39618 55310
rect 35074 55246 35086 55298
rect 35138 55246 35150 55298
rect 35410 55246 35422 55298
rect 35474 55246 35486 55298
rect 37202 55246 37214 55298
rect 37266 55246 37278 55298
rect 38994 55246 39006 55298
rect 39058 55246 39070 55298
rect 40226 55246 40238 55298
rect 40290 55246 40302 55298
rect 48738 55246 48750 55298
rect 48802 55246 48814 55298
rect 51762 55246 51774 55298
rect 51826 55246 51838 55298
rect 52994 55246 53006 55298
rect 53058 55246 53070 55298
rect 34078 55234 34130 55246
rect 36990 55234 37042 55246
rect 39566 55234 39618 55246
rect 19630 55186 19682 55198
rect 19630 55122 19682 55134
rect 19966 55186 20018 55198
rect 19966 55122 20018 55134
rect 20190 55186 20242 55198
rect 25678 55186 25730 55198
rect 24882 55134 24894 55186
rect 24946 55134 24958 55186
rect 20190 55122 20242 55134
rect 25678 55122 25730 55134
rect 26462 55186 26514 55198
rect 26462 55122 26514 55134
rect 27806 55186 27858 55198
rect 27806 55122 27858 55134
rect 30830 55186 30882 55198
rect 37774 55186 37826 55198
rect 32946 55134 32958 55186
rect 33010 55134 33022 55186
rect 34514 55134 34526 55186
rect 34578 55134 34590 55186
rect 30830 55122 30882 55134
rect 37774 55122 37826 55134
rect 41022 55186 41074 55198
rect 41022 55122 41074 55134
rect 42478 55186 42530 55198
rect 42478 55122 42530 55134
rect 44830 55186 44882 55198
rect 44830 55122 44882 55134
rect 45390 55186 45442 55198
rect 45390 55122 45442 55134
rect 45502 55186 45554 55198
rect 45502 55122 45554 55134
rect 45726 55186 45778 55198
rect 45726 55122 45778 55134
rect 46846 55186 46898 55198
rect 46846 55122 46898 55134
rect 46958 55186 47010 55198
rect 46958 55122 47010 55134
rect 47070 55186 47122 55198
rect 47854 55186 47906 55198
rect 47506 55134 47518 55186
rect 47570 55134 47582 55186
rect 47070 55122 47122 55134
rect 47854 55122 47906 55134
rect 57710 55186 57762 55198
rect 57710 55122 57762 55134
rect 18734 55074 18786 55086
rect 18734 55010 18786 55022
rect 19182 55074 19234 55086
rect 19182 55010 19234 55022
rect 19854 55074 19906 55086
rect 19854 55010 19906 55022
rect 20862 55074 20914 55086
rect 20862 55010 20914 55022
rect 21310 55074 21362 55086
rect 22206 55074 22258 55086
rect 21634 55022 21646 55074
rect 21698 55022 21710 55074
rect 21310 55010 21362 55022
rect 22206 55010 22258 55022
rect 22430 55074 22482 55086
rect 25790 55074 25842 55086
rect 22754 55022 22766 55074
rect 22818 55022 22830 55074
rect 22430 55010 22482 55022
rect 25790 55010 25842 55022
rect 26014 55074 26066 55086
rect 26014 55010 26066 55022
rect 26574 55074 26626 55086
rect 26574 55010 26626 55022
rect 26798 55074 26850 55086
rect 26798 55010 26850 55022
rect 27470 55074 27522 55086
rect 27470 55010 27522 55022
rect 27918 55074 27970 55086
rect 27918 55010 27970 55022
rect 28030 55074 28082 55086
rect 28030 55010 28082 55022
rect 28590 55074 28642 55086
rect 30494 55074 30546 55086
rect 42030 55074 42082 55086
rect 30146 55022 30158 55074
rect 30210 55022 30222 55074
rect 31154 55022 31166 55074
rect 31218 55022 31230 55074
rect 35522 55022 35534 55074
rect 35586 55022 35598 55074
rect 28590 55010 28642 55022
rect 30494 55010 30546 55022
rect 42030 55010 42082 55022
rect 42142 55074 42194 55086
rect 42142 55010 42194 55022
rect 42254 55074 42306 55086
rect 42254 55010 42306 55022
rect 44942 55074 44994 55086
rect 44942 55010 44994 55022
rect 45166 55074 45218 55086
rect 45166 55010 45218 55022
rect 48078 55074 48130 55086
rect 48078 55010 48130 55022
rect 51550 55074 51602 55086
rect 51550 55010 51602 55022
rect 58158 55074 58210 55086
rect 58158 55010 58210 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 45054 54738 45106 54750
rect 27234 54686 27246 54738
rect 27298 54686 27310 54738
rect 45054 54674 45106 54686
rect 47406 54738 47458 54750
rect 47406 54674 47458 54686
rect 52334 54738 52386 54750
rect 52334 54674 52386 54686
rect 1710 54626 1762 54638
rect 33182 54626 33234 54638
rect 44718 54626 44770 54638
rect 19394 54574 19406 54626
rect 19458 54574 19470 54626
rect 21298 54574 21310 54626
rect 21362 54574 21374 54626
rect 26338 54574 26350 54626
rect 26402 54574 26414 54626
rect 29362 54574 29374 54626
rect 29426 54574 29438 54626
rect 34178 54574 34190 54626
rect 34242 54574 34254 54626
rect 1710 54562 1762 54574
rect 33182 54562 33234 54574
rect 44718 54562 44770 54574
rect 44830 54626 44882 54638
rect 44830 54562 44882 54574
rect 46846 54626 46898 54638
rect 46846 54562 46898 54574
rect 49086 54626 49138 54638
rect 49086 54562 49138 54574
rect 49310 54626 49362 54638
rect 49310 54562 49362 54574
rect 50878 54626 50930 54638
rect 50878 54562 50930 54574
rect 22206 54514 22258 54526
rect 18610 54462 18622 54514
rect 18674 54462 18686 54514
rect 20402 54462 20414 54514
rect 20466 54462 20478 54514
rect 21186 54462 21198 54514
rect 21250 54462 21262 54514
rect 22206 54450 22258 54462
rect 22430 54514 22482 54526
rect 22430 54450 22482 54462
rect 23326 54514 23378 54526
rect 23326 54450 23378 54462
rect 23662 54514 23714 54526
rect 28142 54514 28194 54526
rect 42254 54514 42306 54526
rect 44382 54514 44434 54526
rect 47070 54514 47122 54526
rect 25890 54462 25902 54514
rect 25954 54462 25966 54514
rect 26786 54462 26798 54514
rect 26850 54462 26862 54514
rect 27122 54462 27134 54514
rect 27186 54462 27198 54514
rect 28466 54462 28478 54514
rect 28530 54462 28542 54514
rect 29026 54462 29038 54514
rect 29090 54462 29102 54514
rect 30594 54462 30606 54514
rect 30658 54462 30670 54514
rect 31938 54462 31950 54514
rect 32002 54462 32014 54514
rect 34066 54462 34078 54514
rect 34130 54462 34142 54514
rect 35634 54462 35646 54514
rect 35698 54462 35710 54514
rect 37202 54462 37214 54514
rect 37266 54462 37278 54514
rect 38098 54462 38110 54514
rect 38162 54462 38174 54514
rect 41570 54462 41582 54514
rect 41634 54462 41646 54514
rect 43474 54462 43486 54514
rect 43538 54462 43550 54514
rect 46386 54462 46398 54514
rect 46450 54462 46462 54514
rect 23662 54450 23714 54462
rect 28142 54450 28194 54462
rect 42254 54450 42306 54462
rect 44382 54450 44434 54462
rect 47070 54450 47122 54462
rect 47518 54514 47570 54526
rect 47518 54450 47570 54462
rect 47630 54514 47682 54526
rect 49970 54462 49982 54514
rect 50034 54462 50046 54514
rect 51538 54462 51550 54514
rect 51602 54462 51614 54514
rect 47630 54450 47682 54462
rect 19070 54402 19122 54414
rect 19070 54338 19122 54350
rect 25678 54402 25730 54414
rect 25678 54338 25730 54350
rect 27918 54402 27970 54414
rect 49198 54402 49250 54414
rect 30146 54350 30158 54402
rect 30210 54350 30222 54402
rect 35186 54350 35198 54402
rect 35250 54350 35262 54402
rect 38434 54350 38446 54402
rect 38498 54350 38510 54402
rect 41346 54350 41358 54402
rect 41410 54350 41422 54402
rect 43810 54350 43822 54402
rect 43874 54350 43886 54402
rect 46162 54350 46174 54402
rect 46226 54350 46238 54402
rect 50194 54350 50206 54402
rect 50258 54350 50270 54402
rect 27918 54338 27970 54350
rect 49198 54338 49250 54350
rect 22094 54290 22146 54302
rect 22094 54226 22146 54238
rect 22654 54290 22706 54302
rect 22654 54226 22706 54238
rect 22766 54290 22818 54302
rect 22766 54226 22818 54238
rect 23438 54290 23490 54302
rect 23438 54226 23490 54238
rect 23774 54290 23826 54302
rect 23774 54226 23826 54238
rect 25566 54290 25618 54302
rect 38658 54238 38670 54290
rect 38722 54238 38734 54290
rect 25566 54226 25618 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 41694 53954 41746 53966
rect 41694 53890 41746 53902
rect 42254 53954 42306 53966
rect 42254 53890 42306 53902
rect 42478 53954 42530 53966
rect 42478 53890 42530 53902
rect 46174 53954 46226 53966
rect 46174 53890 46226 53902
rect 47294 53954 47346 53966
rect 47294 53890 47346 53902
rect 16830 53842 16882 53854
rect 23774 53842 23826 53854
rect 19730 53790 19742 53842
rect 19794 53790 19806 53842
rect 21410 53790 21422 53842
rect 21474 53790 21486 53842
rect 16830 53778 16882 53790
rect 23774 53778 23826 53790
rect 23886 53842 23938 53854
rect 23886 53778 23938 53790
rect 28478 53842 28530 53854
rect 36094 53842 36146 53854
rect 37998 53842 38050 53854
rect 41358 53842 41410 53854
rect 50206 53842 50258 53854
rect 32946 53790 32958 53842
rect 33010 53790 33022 53842
rect 34626 53790 34638 53842
rect 34690 53790 34702 53842
rect 37314 53790 37326 53842
rect 37378 53790 37390 53842
rect 39778 53790 39790 53842
rect 39842 53790 39854 53842
rect 46498 53790 46510 53842
rect 46562 53790 46574 53842
rect 47842 53790 47854 53842
rect 47906 53790 47918 53842
rect 51314 53790 51326 53842
rect 51378 53790 51390 53842
rect 28478 53778 28530 53790
rect 36094 53778 36146 53790
rect 37998 53778 38050 53790
rect 41358 53778 41410 53790
rect 50206 53778 50258 53790
rect 19294 53730 19346 53742
rect 24782 53730 24834 53742
rect 16930 53678 16942 53730
rect 16994 53678 17006 53730
rect 19842 53678 19854 53730
rect 19906 53678 19918 53730
rect 21746 53678 21758 53730
rect 21810 53678 21822 53730
rect 22306 53678 22318 53730
rect 22370 53678 22382 53730
rect 22530 53678 22542 53730
rect 22594 53678 22606 53730
rect 22866 53678 22878 53730
rect 22930 53678 22942 53730
rect 19294 53666 19346 53678
rect 24782 53666 24834 53678
rect 25118 53730 25170 53742
rect 25118 53666 25170 53678
rect 25790 53730 25842 53742
rect 25790 53666 25842 53678
rect 26126 53730 26178 53742
rect 34414 53730 34466 53742
rect 35870 53730 35922 53742
rect 42030 53730 42082 53742
rect 27906 53678 27918 53730
rect 27970 53678 27982 53730
rect 29362 53678 29374 53730
rect 29426 53678 29438 53730
rect 30034 53678 30046 53730
rect 30098 53678 30110 53730
rect 30930 53678 30942 53730
rect 30994 53678 31006 53730
rect 33282 53678 33294 53730
rect 33346 53678 33358 53730
rect 33842 53678 33854 53730
rect 33906 53678 33918 53730
rect 34962 53678 34974 53730
rect 35026 53678 35038 53730
rect 37202 53678 37214 53730
rect 37266 53678 37278 53730
rect 38770 53678 38782 53730
rect 38834 53678 38846 53730
rect 39890 53678 39902 53730
rect 39954 53678 39966 53730
rect 26126 53666 26178 53678
rect 34414 53666 34466 53678
rect 35870 53666 35922 53678
rect 42030 53666 42082 53678
rect 42926 53730 42978 53742
rect 47182 53730 47234 53742
rect 49646 53730 49698 53742
rect 46946 53678 46958 53730
rect 47010 53678 47022 53730
rect 47954 53678 47966 53730
rect 48018 53678 48030 53730
rect 42926 53666 42978 53678
rect 47182 53666 47234 53678
rect 49646 53666 49698 53678
rect 50094 53730 50146 53742
rect 50978 53678 50990 53730
rect 51042 53678 51054 53730
rect 50094 53666 50146 53678
rect 16046 53618 16098 53630
rect 16046 53554 16098 53566
rect 16718 53618 16770 53630
rect 23998 53618 24050 53630
rect 17826 53566 17838 53618
rect 17890 53566 17902 53618
rect 16718 53554 16770 53566
rect 23998 53554 24050 53566
rect 25454 53618 25506 53630
rect 25454 53554 25506 53566
rect 27022 53618 27074 53630
rect 27022 53554 27074 53566
rect 28366 53618 28418 53630
rect 43598 53618 43650 53630
rect 29250 53566 29262 53618
rect 29314 53566 29326 53618
rect 30258 53566 30270 53618
rect 30322 53566 30334 53618
rect 33394 53566 33406 53618
rect 33458 53566 33470 53618
rect 34178 53566 34190 53618
rect 34242 53566 34254 53618
rect 39442 53566 39454 53618
rect 39506 53566 39518 53618
rect 28366 53554 28418 53566
rect 43598 53554 43650 53566
rect 43710 53618 43762 53630
rect 43710 53554 43762 53566
rect 43934 53618 43986 53630
rect 43934 53554 43986 53566
rect 48750 53618 48802 53630
rect 48750 53554 48802 53566
rect 49086 53618 49138 53630
rect 49086 53554 49138 53566
rect 49422 53618 49474 53630
rect 49422 53554 49474 53566
rect 51662 53618 51714 53630
rect 51662 53554 51714 53566
rect 52670 53618 52722 53630
rect 52670 53554 52722 53566
rect 53006 53618 53058 53630
rect 53006 53554 53058 53566
rect 16494 53506 16546 53518
rect 16494 53442 16546 53454
rect 17166 53506 17218 53518
rect 17166 53442 17218 53454
rect 17502 53506 17554 53518
rect 17502 53442 17554 53454
rect 19406 53506 19458 53518
rect 19406 53442 19458 53454
rect 19630 53506 19682 53518
rect 19630 53442 19682 53454
rect 20414 53506 20466 53518
rect 20414 53442 20466 53454
rect 20750 53506 20802 53518
rect 25118 53506 25170 53518
rect 23090 53454 23102 53506
rect 23154 53454 23166 53506
rect 20750 53442 20802 53454
rect 25118 53442 25170 53454
rect 25902 53506 25954 53518
rect 25902 53442 25954 53454
rect 26910 53506 26962 53518
rect 26910 53442 26962 53454
rect 27694 53506 27746 53518
rect 27694 53442 27746 53454
rect 28142 53506 28194 53518
rect 28142 53442 28194 53454
rect 31502 53506 31554 53518
rect 41582 53506 41634 53518
rect 36418 53454 36430 53506
rect 36482 53454 36494 53506
rect 31502 53442 31554 53454
rect 41582 53442 41634 53454
rect 46398 53506 46450 53518
rect 46398 53442 46450 53454
rect 50318 53506 50370 53518
rect 50318 53442 50370 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 20414 53170 20466 53182
rect 20414 53106 20466 53118
rect 22766 53170 22818 53182
rect 22766 53106 22818 53118
rect 23326 53170 23378 53182
rect 23326 53106 23378 53118
rect 27806 53170 27858 53182
rect 27806 53106 27858 53118
rect 28814 53170 28866 53182
rect 28814 53106 28866 53118
rect 30830 53170 30882 53182
rect 30830 53106 30882 53118
rect 33630 53170 33682 53182
rect 33630 53106 33682 53118
rect 38894 53170 38946 53182
rect 38894 53106 38946 53118
rect 39006 53170 39058 53182
rect 39006 53106 39058 53118
rect 17502 53058 17554 53070
rect 18846 53058 18898 53070
rect 16594 53006 16606 53058
rect 16658 53006 16670 53058
rect 18610 53006 18622 53058
rect 18674 53006 18686 53058
rect 17502 52994 17554 53006
rect 18846 52994 18898 53006
rect 19630 53058 19682 53070
rect 19630 52994 19682 53006
rect 20638 53058 20690 53070
rect 20638 52994 20690 53006
rect 20750 53058 20802 53070
rect 31278 53058 31330 53070
rect 28130 53006 28142 53058
rect 28194 53006 28206 53058
rect 20750 52994 20802 53006
rect 31278 52994 31330 53006
rect 38782 53058 38834 53070
rect 38782 52994 38834 53006
rect 50654 53058 50706 53070
rect 50654 52994 50706 53006
rect 58158 53058 58210 53070
rect 58158 52994 58210 53006
rect 17278 52946 17330 52958
rect 16706 52894 16718 52946
rect 16770 52894 16782 52946
rect 17278 52882 17330 52894
rect 17614 52946 17666 52958
rect 17614 52882 17666 52894
rect 18398 52946 18450 52958
rect 18398 52882 18450 52894
rect 18510 52946 18562 52958
rect 18510 52882 18562 52894
rect 19294 52946 19346 52958
rect 19294 52882 19346 52894
rect 22094 52946 22146 52958
rect 22094 52882 22146 52894
rect 22542 52946 22594 52958
rect 22542 52882 22594 52894
rect 31054 52946 31106 52958
rect 31054 52882 31106 52894
rect 31950 52946 32002 52958
rect 31950 52882 32002 52894
rect 33406 52946 33458 52958
rect 33406 52882 33458 52894
rect 33742 52946 33794 52958
rect 36766 52946 36818 52958
rect 34178 52894 34190 52946
rect 34242 52894 34254 52946
rect 34738 52894 34750 52946
rect 34802 52894 34814 52946
rect 33742 52882 33794 52894
rect 36766 52882 36818 52894
rect 47182 52946 47234 52958
rect 47182 52882 47234 52894
rect 47406 52946 47458 52958
rect 50978 52894 50990 52946
rect 51042 52894 51054 52946
rect 51762 52894 51774 52946
rect 51826 52894 51838 52946
rect 47406 52882 47458 52894
rect 21198 52834 21250 52846
rect 21198 52770 21250 52782
rect 22318 52834 22370 52846
rect 24558 52834 24610 52846
rect 22642 52782 22654 52834
rect 22706 52782 22718 52834
rect 22318 52770 22370 52782
rect 24558 52770 24610 52782
rect 26462 52834 26514 52846
rect 26462 52770 26514 52782
rect 29262 52834 29314 52846
rect 29262 52770 29314 52782
rect 30942 52834 30994 52846
rect 30942 52770 30994 52782
rect 31726 52834 31778 52846
rect 31726 52770 31778 52782
rect 32286 52834 32338 52846
rect 34626 52782 34638 52834
rect 34690 52782 34702 52834
rect 36306 52782 36318 52834
rect 36370 52782 36382 52834
rect 50866 52782 50878 52834
rect 50930 52782 50942 52834
rect 51650 52782 51662 52834
rect 51714 52782 51726 52834
rect 32286 52770 32338 52782
rect 15598 52722 15650 52734
rect 15598 52658 15650 52670
rect 15934 52722 15986 52734
rect 15934 52658 15986 52670
rect 19182 52722 19234 52734
rect 19182 52658 19234 52670
rect 19742 52722 19794 52734
rect 19742 52658 19794 52670
rect 19966 52722 20018 52734
rect 19966 52658 20018 52670
rect 20078 52722 20130 52734
rect 20078 52658 20130 52670
rect 21870 52722 21922 52734
rect 47630 52722 47682 52734
rect 35074 52670 35086 52722
rect 35138 52670 35150 52722
rect 21870 52658 21922 52670
rect 47630 52658 47682 52670
rect 48078 52722 48130 52734
rect 48078 52658 48130 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 22990 52386 23042 52398
rect 22990 52322 23042 52334
rect 23438 52386 23490 52398
rect 23438 52322 23490 52334
rect 31278 52386 31330 52398
rect 47966 52386 48018 52398
rect 43586 52334 43598 52386
rect 43650 52334 43662 52386
rect 31278 52322 31330 52334
rect 47966 52322 48018 52334
rect 15822 52274 15874 52286
rect 15822 52210 15874 52222
rect 19070 52274 19122 52286
rect 21422 52274 21474 52286
rect 19618 52222 19630 52274
rect 19682 52222 19694 52274
rect 19070 52210 19122 52222
rect 21422 52210 21474 52222
rect 25342 52274 25394 52286
rect 25342 52210 25394 52222
rect 27470 52274 27522 52286
rect 27470 52210 27522 52222
rect 34190 52274 34242 52286
rect 34190 52210 34242 52222
rect 40014 52274 40066 52286
rect 40014 52210 40066 52222
rect 40910 52274 40962 52286
rect 51326 52274 51378 52286
rect 43250 52222 43262 52274
rect 43314 52222 43326 52274
rect 40910 52210 40962 52222
rect 51326 52210 51378 52222
rect 51774 52274 51826 52286
rect 51774 52210 51826 52222
rect 16382 52162 16434 52174
rect 16382 52098 16434 52110
rect 16942 52162 16994 52174
rect 16942 52098 16994 52110
rect 19406 52162 19458 52174
rect 19406 52098 19458 52110
rect 20862 52162 20914 52174
rect 23662 52162 23714 52174
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 22082 52110 22094 52162
rect 22146 52110 22158 52162
rect 22754 52110 22766 52162
rect 22818 52110 22830 52162
rect 20862 52098 20914 52110
rect 23662 52098 23714 52110
rect 23998 52162 24050 52174
rect 30494 52162 30546 52174
rect 24546 52110 24558 52162
rect 24610 52110 24622 52162
rect 25554 52110 25566 52162
rect 25618 52110 25630 52162
rect 26898 52110 26910 52162
rect 26962 52110 26974 52162
rect 27682 52110 27694 52162
rect 27746 52110 27758 52162
rect 28690 52159 28702 52162
rect 28481 52113 28702 52159
rect 23998 52098 24050 52110
rect 20526 52050 20578 52062
rect 20526 51986 20578 51998
rect 20638 52050 20690 52062
rect 24994 51998 25006 52050
rect 25058 51998 25070 52050
rect 25330 51998 25342 52050
rect 25394 51998 25406 52050
rect 27122 51998 27134 52050
rect 27186 51998 27198 52050
rect 28354 51998 28366 52050
rect 28418 52047 28430 52050
rect 28481 52047 28527 52113
rect 28690 52110 28702 52113
rect 28754 52110 28766 52162
rect 30494 52098 30546 52110
rect 34078 52162 34130 52174
rect 34078 52098 34130 52110
rect 34302 52162 34354 52174
rect 34302 52098 34354 52110
rect 34638 52162 34690 52174
rect 39118 52162 39170 52174
rect 38434 52110 38446 52162
rect 38498 52110 38510 52162
rect 34638 52098 34690 52110
rect 39118 52098 39170 52110
rect 40574 52162 40626 52174
rect 40574 52098 40626 52110
rect 42030 52162 42082 52174
rect 51438 52162 51490 52174
rect 42242 52110 42254 52162
rect 42306 52110 42318 52162
rect 43138 52110 43150 52162
rect 43202 52110 43214 52162
rect 43474 52110 43486 52162
rect 43538 52110 43550 52162
rect 42030 52098 42082 52110
rect 51438 52098 51490 52110
rect 28418 52001 28527 52047
rect 31166 52050 31218 52062
rect 28418 51998 28430 52001
rect 20638 51986 20690 51998
rect 31166 51986 31218 51998
rect 31278 52050 31330 52062
rect 45726 52050 45778 52062
rect 38546 51998 38558 52050
rect 38610 51998 38622 52050
rect 31278 51986 31330 51998
rect 45726 51986 45778 51998
rect 47630 52050 47682 52062
rect 47630 51986 47682 51998
rect 47854 52050 47906 52062
rect 47854 51986 47906 51998
rect 15486 51938 15538 51950
rect 15486 51874 15538 51886
rect 15710 51938 15762 51950
rect 15710 51874 15762 51886
rect 15934 51938 15986 51950
rect 15934 51874 15986 51886
rect 23886 51938 23938 51950
rect 23886 51874 23938 51886
rect 24110 51938 24162 51950
rect 29262 51938 29314 51950
rect 39454 51938 39506 51950
rect 27234 51886 27246 51938
rect 27298 51886 27310 51938
rect 30818 51886 30830 51938
rect 30882 51886 30894 51938
rect 24110 51874 24162 51886
rect 29262 51874 29314 51886
rect 39454 51874 39506 51886
rect 39902 51938 39954 51950
rect 39902 51874 39954 51886
rect 40126 51938 40178 51950
rect 40126 51874 40178 51886
rect 40798 51938 40850 51950
rect 40798 51874 40850 51886
rect 41022 51938 41074 51950
rect 41022 51874 41074 51886
rect 41246 51938 41298 51950
rect 41246 51874 41298 51886
rect 45838 51938 45890 51950
rect 45838 51874 45890 51886
rect 46062 51938 46114 51950
rect 46062 51874 46114 51886
rect 50990 51938 51042 51950
rect 50990 51874 51042 51886
rect 51214 51938 51266 51950
rect 51214 51874 51266 51886
rect 51886 51938 51938 51950
rect 51886 51874 51938 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 23886 51602 23938 51614
rect 22978 51550 22990 51602
rect 23042 51550 23054 51602
rect 23886 51538 23938 51550
rect 24558 51602 24610 51614
rect 24558 51538 24610 51550
rect 25678 51602 25730 51614
rect 25678 51538 25730 51550
rect 39454 51602 39506 51614
rect 39454 51538 39506 51550
rect 41022 51602 41074 51614
rect 41022 51538 41074 51550
rect 47294 51602 47346 51614
rect 51650 51550 51662 51602
rect 51714 51550 51726 51602
rect 47294 51538 47346 51550
rect 16494 51490 16546 51502
rect 23662 51490 23714 51502
rect 19170 51438 19182 51490
rect 19234 51438 19246 51490
rect 23202 51438 23214 51490
rect 23266 51438 23278 51490
rect 16494 51426 16546 51438
rect 23662 51426 23714 51438
rect 28366 51490 28418 51502
rect 28366 51426 28418 51438
rect 28478 51490 28530 51502
rect 28478 51426 28530 51438
rect 36990 51490 37042 51502
rect 36990 51426 37042 51438
rect 37550 51490 37602 51502
rect 41134 51490 41186 51502
rect 38322 51438 38334 51490
rect 38386 51438 38398 51490
rect 38770 51438 38782 51490
rect 38834 51438 38846 51490
rect 37550 51426 37602 51438
rect 41134 51426 41186 51438
rect 42702 51490 42754 51502
rect 42702 51426 42754 51438
rect 46174 51490 46226 51502
rect 46174 51426 46226 51438
rect 47406 51490 47458 51502
rect 53902 51490 53954 51502
rect 51090 51438 51102 51490
rect 51154 51438 51166 51490
rect 47406 51426 47458 51438
rect 53902 51426 53954 51438
rect 58158 51490 58210 51502
rect 58158 51426 58210 51438
rect 15486 51378 15538 51390
rect 16718 51378 16770 51390
rect 24110 51378 24162 51390
rect 15138 51326 15150 51378
rect 15202 51326 15214 51378
rect 15922 51326 15934 51378
rect 15986 51326 15998 51378
rect 16258 51326 16270 51378
rect 16322 51326 16334 51378
rect 19058 51326 19070 51378
rect 19122 51326 19134 51378
rect 20962 51326 20974 51378
rect 21026 51326 21038 51378
rect 22530 51326 22542 51378
rect 22594 51326 22606 51378
rect 15486 51314 15538 51326
rect 16718 51314 16770 51326
rect 24110 51314 24162 51326
rect 25118 51378 25170 51390
rect 25118 51314 25170 51326
rect 25566 51378 25618 51390
rect 25566 51314 25618 51326
rect 25790 51378 25842 51390
rect 25790 51314 25842 51326
rect 26462 51378 26514 51390
rect 27806 51378 27858 51390
rect 27234 51326 27246 51378
rect 27298 51326 27310 51378
rect 26462 51314 26514 51326
rect 27806 51314 27858 51326
rect 28142 51378 28194 51390
rect 29262 51378 29314 51390
rect 28914 51326 28926 51378
rect 28978 51326 28990 51378
rect 28142 51314 28194 51326
rect 29262 51314 29314 51326
rect 30606 51378 30658 51390
rect 30606 51314 30658 51326
rect 30830 51378 30882 51390
rect 30830 51314 30882 51326
rect 31054 51378 31106 51390
rect 31054 51314 31106 51326
rect 31278 51378 31330 51390
rect 36094 51378 36146 51390
rect 39118 51378 39170 51390
rect 46958 51378 47010 51390
rect 34290 51326 34302 51378
rect 34354 51326 34366 51378
rect 36418 51326 36430 51378
rect 36482 51326 36494 51378
rect 37874 51326 37886 51378
rect 37938 51326 37950 51378
rect 42018 51326 42030 51378
rect 42082 51326 42094 51378
rect 43362 51326 43374 51378
rect 43426 51326 43438 51378
rect 45714 51326 45726 51378
rect 45778 51326 45790 51378
rect 31278 51314 31330 51326
rect 36094 51314 36146 51326
rect 39118 51314 39170 51326
rect 46958 51314 47010 51326
rect 47070 51378 47122 51390
rect 53230 51378 53282 51390
rect 50866 51326 50878 51378
rect 50930 51326 50942 51378
rect 51538 51326 51550 51378
rect 51602 51326 51614 51378
rect 52770 51326 52782 51378
rect 52834 51326 52846 51378
rect 47070 51314 47122 51326
rect 53230 51314 53282 51326
rect 53566 51378 53618 51390
rect 53566 51314 53618 51326
rect 15598 51266 15650 51278
rect 17502 51266 17554 51278
rect 16370 51214 16382 51266
rect 16434 51214 16446 51266
rect 15598 51202 15650 51214
rect 17502 51202 17554 51214
rect 18398 51266 18450 51278
rect 18398 51202 18450 51214
rect 18734 51266 18786 51278
rect 18734 51202 18786 51214
rect 23998 51266 24050 51278
rect 28254 51266 28306 51278
rect 26898 51214 26910 51266
rect 26962 51214 26974 51266
rect 23998 51202 24050 51214
rect 28254 51202 28306 51214
rect 29822 51266 29874 51278
rect 29822 51202 29874 51214
rect 31166 51266 31218 51278
rect 44046 51266 44098 51278
rect 34066 51214 34078 51266
rect 34130 51214 34142 51266
rect 42242 51214 42254 51266
rect 42306 51214 42318 51266
rect 43250 51214 43262 51266
rect 43314 51214 43326 51266
rect 45490 51214 45502 51266
rect 45554 51214 45566 51266
rect 52322 51214 52334 51266
rect 52386 51214 52398 51266
rect 31166 51202 31218 51214
rect 44046 51202 44098 51214
rect 37886 51154 37938 51166
rect 24322 51102 24334 51154
rect 24386 51151 24398 51154
rect 24770 51151 24782 51154
rect 24386 51105 24782 51151
rect 24386 51102 24398 51105
rect 24770 51102 24782 51105
rect 24834 51102 24846 51154
rect 34738 51102 34750 51154
rect 34802 51102 34814 51154
rect 37886 51090 37938 51102
rect 40910 51154 40962 51166
rect 40910 51090 40962 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 17726 50818 17778 50830
rect 15474 50766 15486 50818
rect 15538 50815 15550 50818
rect 16370 50815 16382 50818
rect 15538 50769 16382 50815
rect 15538 50766 15550 50769
rect 16370 50766 16382 50769
rect 16434 50766 16446 50818
rect 17726 50754 17778 50766
rect 18062 50818 18114 50830
rect 18062 50754 18114 50766
rect 19518 50818 19570 50830
rect 19518 50754 19570 50766
rect 25342 50818 25394 50830
rect 25342 50754 25394 50766
rect 34862 50818 34914 50830
rect 34862 50754 34914 50766
rect 42142 50818 42194 50830
rect 42142 50754 42194 50766
rect 42478 50818 42530 50830
rect 52782 50818 52834 50830
rect 47394 50766 47406 50818
rect 47458 50766 47470 50818
rect 42478 50754 42530 50766
rect 52782 50754 52834 50766
rect 57934 50818 57986 50830
rect 57934 50754 57986 50766
rect 12910 50706 12962 50718
rect 17390 50706 17442 50718
rect 15138 50654 15150 50706
rect 15202 50654 15214 50706
rect 12910 50642 12962 50654
rect 17390 50642 17442 50654
rect 20190 50706 20242 50718
rect 20190 50642 20242 50654
rect 22542 50706 22594 50718
rect 22542 50642 22594 50654
rect 23886 50706 23938 50718
rect 23886 50642 23938 50654
rect 27582 50706 27634 50718
rect 27582 50642 27634 50654
rect 39230 50706 39282 50718
rect 44930 50654 44942 50706
rect 44994 50654 45006 50706
rect 39230 50642 39282 50654
rect 13470 50594 13522 50606
rect 13470 50530 13522 50542
rect 14142 50594 14194 50606
rect 14142 50530 14194 50542
rect 18846 50594 18898 50606
rect 18846 50530 18898 50542
rect 22094 50594 22146 50606
rect 22094 50530 22146 50542
rect 22318 50594 22370 50606
rect 25566 50594 25618 50606
rect 29486 50594 29538 50606
rect 25218 50542 25230 50594
rect 25282 50542 25294 50594
rect 29138 50542 29150 50594
rect 29202 50542 29214 50594
rect 22318 50530 22370 50542
rect 25566 50530 25618 50542
rect 29486 50530 29538 50542
rect 31166 50594 31218 50606
rect 31166 50530 31218 50542
rect 33294 50594 33346 50606
rect 34526 50594 34578 50606
rect 33954 50542 33966 50594
rect 34018 50542 34030 50594
rect 33294 50530 33346 50542
rect 34526 50530 34578 50542
rect 38782 50594 38834 50606
rect 38782 50530 38834 50542
rect 39342 50594 39394 50606
rect 44046 50594 44098 50606
rect 46846 50594 46898 50606
rect 51662 50594 51714 50606
rect 42466 50542 42478 50594
rect 42530 50542 42542 50594
rect 45154 50542 45166 50594
rect 45218 50542 45230 50594
rect 46610 50542 46622 50594
rect 46674 50542 46686 50594
rect 47730 50542 47742 50594
rect 47794 50542 47806 50594
rect 48626 50542 48638 50594
rect 48690 50542 48702 50594
rect 50418 50542 50430 50594
rect 50482 50542 50494 50594
rect 39342 50530 39394 50542
rect 44046 50530 44098 50542
rect 46846 50530 46898 50542
rect 51662 50530 51714 50542
rect 52894 50594 52946 50606
rect 55570 50542 55582 50594
rect 55634 50542 55646 50594
rect 52894 50530 52946 50542
rect 14590 50482 14642 50494
rect 14590 50418 14642 50430
rect 14814 50482 14866 50494
rect 14814 50418 14866 50430
rect 15038 50482 15090 50494
rect 15038 50418 15090 50430
rect 15262 50482 15314 50494
rect 18622 50482 18674 50494
rect 16930 50430 16942 50482
rect 16994 50430 17006 50482
rect 15262 50418 15314 50430
rect 18622 50418 18674 50430
rect 19406 50482 19458 50494
rect 19406 50418 19458 50430
rect 19518 50482 19570 50494
rect 19518 50418 19570 50430
rect 20526 50482 20578 50494
rect 20526 50418 20578 50430
rect 20638 50482 20690 50494
rect 20638 50418 20690 50430
rect 20862 50482 20914 50494
rect 20862 50418 20914 50430
rect 22654 50482 22706 50494
rect 22654 50418 22706 50430
rect 22990 50482 23042 50494
rect 22990 50418 23042 50430
rect 23102 50482 23154 50494
rect 23102 50418 23154 50430
rect 23774 50482 23826 50494
rect 23774 50418 23826 50430
rect 25006 50482 25058 50494
rect 25006 50418 25058 50430
rect 26462 50482 26514 50494
rect 26462 50418 26514 50430
rect 27694 50482 27746 50494
rect 27694 50418 27746 50430
rect 28142 50482 28194 50494
rect 28142 50418 28194 50430
rect 30382 50482 30434 50494
rect 30382 50418 30434 50430
rect 31054 50482 31106 50494
rect 31054 50418 31106 50430
rect 31502 50482 31554 50494
rect 31502 50418 31554 50430
rect 31726 50482 31778 50494
rect 31726 50418 31778 50430
rect 31838 50482 31890 50494
rect 31838 50418 31890 50430
rect 32958 50482 33010 50494
rect 32958 50418 33010 50430
rect 33070 50482 33122 50494
rect 39006 50482 39058 50494
rect 33842 50430 33854 50482
rect 33906 50430 33918 50482
rect 33070 50418 33122 50430
rect 39006 50418 39058 50430
rect 39902 50482 39954 50494
rect 39902 50418 39954 50430
rect 44158 50482 44210 50494
rect 44158 50418 44210 50430
rect 44382 50482 44434 50494
rect 44382 50418 44434 50430
rect 45838 50482 45890 50494
rect 45838 50418 45890 50430
rect 46958 50482 47010 50494
rect 52782 50482 52834 50494
rect 48066 50430 48078 50482
rect 48130 50430 48142 50482
rect 50754 50430 50766 50482
rect 50818 50430 50830 50482
rect 51090 50430 51102 50482
rect 51154 50430 51166 50482
rect 46958 50418 47010 50430
rect 52782 50418 52834 50430
rect 13582 50370 13634 50382
rect 13582 50306 13634 50318
rect 13694 50370 13746 50382
rect 13694 50306 13746 50318
rect 15710 50370 15762 50382
rect 15710 50306 15762 50318
rect 16382 50370 16434 50382
rect 16382 50306 16434 50318
rect 16606 50370 16658 50382
rect 16606 50306 16658 50318
rect 17950 50370 18002 50382
rect 17950 50306 18002 50318
rect 18958 50370 19010 50382
rect 18958 50306 19010 50318
rect 19182 50370 19234 50382
rect 19182 50306 19234 50318
rect 21422 50370 21474 50382
rect 21422 50306 21474 50318
rect 23326 50370 23378 50382
rect 23326 50306 23378 50318
rect 23998 50370 24050 50382
rect 23998 50306 24050 50318
rect 28702 50370 28754 50382
rect 28702 50306 28754 50318
rect 29598 50370 29650 50382
rect 29598 50306 29650 50318
rect 29710 50370 29762 50382
rect 48626 50318 48638 50370
rect 48690 50318 48702 50370
rect 29710 50306 29762 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 19294 50034 19346 50046
rect 29822 50034 29874 50046
rect 21074 49982 21086 50034
rect 21138 49982 21150 50034
rect 27010 49982 27022 50034
rect 27074 49982 27086 50034
rect 19294 49970 19346 49982
rect 29822 49970 29874 49982
rect 30606 50034 30658 50046
rect 30606 49970 30658 49982
rect 34190 50034 34242 50046
rect 34190 49970 34242 49982
rect 35422 50034 35474 50046
rect 35422 49970 35474 49982
rect 38110 50034 38162 50046
rect 38110 49970 38162 49982
rect 47518 50034 47570 50046
rect 50418 49982 50430 50034
rect 50482 49982 50494 50034
rect 47518 49970 47570 49982
rect 12462 49922 12514 49934
rect 12462 49858 12514 49870
rect 16270 49922 16322 49934
rect 16270 49858 16322 49870
rect 16382 49922 16434 49934
rect 16382 49858 16434 49870
rect 17838 49922 17890 49934
rect 17838 49858 17890 49870
rect 18398 49922 18450 49934
rect 18398 49858 18450 49870
rect 19630 49922 19682 49934
rect 21198 49922 21250 49934
rect 20402 49870 20414 49922
rect 20466 49870 20478 49922
rect 19630 49858 19682 49870
rect 21198 49858 21250 49870
rect 24110 49922 24162 49934
rect 30046 49922 30098 49934
rect 25330 49870 25342 49922
rect 25394 49870 25406 49922
rect 24110 49858 24162 49870
rect 30046 49858 30098 49870
rect 35534 49922 35586 49934
rect 43038 49922 43090 49934
rect 36866 49870 36878 49922
rect 36930 49870 36942 49922
rect 39890 49870 39902 49922
rect 39954 49870 39966 49922
rect 35534 49858 35586 49870
rect 43038 49858 43090 49870
rect 43150 49922 43202 49934
rect 43150 49858 43202 49870
rect 45054 49922 45106 49934
rect 45054 49858 45106 49870
rect 46846 49922 46898 49934
rect 46846 49858 46898 49870
rect 47854 49922 47906 49934
rect 47854 49858 47906 49870
rect 58158 49922 58210 49934
rect 58158 49858 58210 49870
rect 16046 49810 16098 49822
rect 17502 49810 17554 49822
rect 13122 49758 13134 49810
rect 13186 49758 13198 49810
rect 13794 49758 13806 49810
rect 13858 49758 13870 49810
rect 16706 49758 16718 49810
rect 16770 49758 16782 49810
rect 16046 49746 16098 49758
rect 17502 49746 17554 49758
rect 18958 49810 19010 49822
rect 18958 49746 19010 49758
rect 19406 49810 19458 49822
rect 26686 49810 26738 49822
rect 20178 49758 20190 49810
rect 20242 49758 20254 49810
rect 21410 49758 21422 49810
rect 21474 49758 21486 49810
rect 21858 49758 21870 49810
rect 21922 49758 21934 49810
rect 22418 49758 22430 49810
rect 22482 49758 22494 49810
rect 23202 49758 23214 49810
rect 23266 49758 23278 49810
rect 25218 49758 25230 49810
rect 25282 49758 25294 49810
rect 26114 49758 26126 49810
rect 26178 49758 26190 49810
rect 19406 49746 19458 49758
rect 26686 49746 26738 49758
rect 28030 49810 28082 49822
rect 30718 49810 30770 49822
rect 29586 49758 29598 49810
rect 29650 49758 29662 49810
rect 30258 49758 30270 49810
rect 30322 49758 30334 49810
rect 28030 49746 28082 49758
rect 30718 49746 30770 49758
rect 30830 49810 30882 49822
rect 37438 49810 37490 49822
rect 31154 49758 31166 49810
rect 31218 49758 31230 49810
rect 34402 49758 34414 49810
rect 34466 49758 34478 49810
rect 35746 49758 35758 49810
rect 35810 49758 35822 49810
rect 36530 49758 36542 49810
rect 36594 49758 36606 49810
rect 30830 49746 30882 49758
rect 37438 49746 37490 49758
rect 37886 49810 37938 49822
rect 37886 49746 37938 49758
rect 39566 49810 39618 49822
rect 39566 49746 39618 49758
rect 43374 49810 43426 49822
rect 47182 49810 47234 49822
rect 45378 49758 45390 49810
rect 45442 49758 45454 49810
rect 45938 49758 45950 49810
rect 46002 49758 46014 49810
rect 43374 49746 43426 49758
rect 47182 49746 47234 49758
rect 47630 49810 47682 49822
rect 47630 49746 47682 49758
rect 49870 49810 49922 49822
rect 49870 49746 49922 49758
rect 11230 49698 11282 49710
rect 11230 49634 11282 49646
rect 11678 49698 11730 49710
rect 11678 49634 11730 49646
rect 12126 49698 12178 49710
rect 14702 49698 14754 49710
rect 13458 49646 13470 49698
rect 13522 49646 13534 49698
rect 12126 49634 12178 49646
rect 14702 49634 14754 49646
rect 15710 49698 15762 49710
rect 23550 49698 23602 49710
rect 24670 49698 24722 49710
rect 28590 49698 28642 49710
rect 16818 49646 16830 49698
rect 16882 49646 16894 49698
rect 24210 49646 24222 49698
rect 24274 49646 24286 49698
rect 25442 49646 25454 49698
rect 25506 49646 25518 49698
rect 15710 49634 15762 49646
rect 23550 49634 23602 49646
rect 24670 49634 24722 49646
rect 28590 49634 28642 49646
rect 29262 49698 29314 49710
rect 37998 49698 38050 49710
rect 50094 49698 50146 49710
rect 30034 49646 30046 49698
rect 30098 49646 30110 49698
rect 36418 49646 36430 49698
rect 36482 49646 36494 49698
rect 46050 49646 46062 49698
rect 46114 49646 46126 49698
rect 29262 49634 29314 49646
rect 37998 49634 38050 49646
rect 50094 49634 50146 49646
rect 12014 49586 12066 49598
rect 11106 49534 11118 49586
rect 11170 49583 11182 49586
rect 11666 49583 11678 49586
rect 11170 49537 11678 49583
rect 11170 49534 11182 49537
rect 11666 49534 11678 49537
rect 11730 49534 11742 49586
rect 12014 49522 12066 49534
rect 12350 49586 12402 49598
rect 12350 49522 12402 49534
rect 14030 49586 14082 49598
rect 14030 49522 14082 49534
rect 22990 49586 23042 49598
rect 22990 49522 23042 49534
rect 23886 49586 23938 49598
rect 23886 49522 23938 49534
rect 34078 49586 34130 49598
rect 34078 49522 34130 49534
rect 35422 49586 35474 49598
rect 35422 49522 35474 49534
rect 45390 49586 45442 49598
rect 45390 49522 45442 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 44270 49250 44322 49262
rect 19730 49198 19742 49250
rect 19794 49198 19806 49250
rect 35858 49198 35870 49250
rect 35922 49198 35934 49250
rect 44270 49186 44322 49198
rect 47854 49250 47906 49262
rect 50990 49250 51042 49262
rect 49746 49198 49758 49250
rect 49810 49198 49822 49250
rect 47854 49186 47906 49198
rect 50990 49186 51042 49198
rect 14590 49138 14642 49150
rect 20750 49138 20802 49150
rect 13570 49086 13582 49138
rect 13634 49086 13646 49138
rect 17826 49086 17838 49138
rect 17890 49086 17902 49138
rect 19282 49086 19294 49138
rect 19346 49086 19358 49138
rect 14590 49074 14642 49086
rect 20750 49074 20802 49086
rect 21758 49138 21810 49150
rect 21758 49074 21810 49086
rect 29262 49138 29314 49150
rect 29262 49074 29314 49086
rect 39006 49138 39058 49150
rect 40238 49138 40290 49150
rect 48974 49138 49026 49150
rect 58158 49138 58210 49150
rect 39554 49086 39566 49138
rect 39618 49086 39630 49138
rect 43586 49086 43598 49138
rect 43650 49086 43662 49138
rect 50082 49086 50094 49138
rect 50146 49086 50158 49138
rect 39006 49074 39058 49086
rect 40238 49074 40290 49086
rect 48974 49074 49026 49086
rect 58158 49074 58210 49086
rect 16606 49026 16658 49038
rect 21646 49026 21698 49038
rect 16146 48974 16158 49026
rect 16210 48974 16222 49026
rect 17154 48974 17166 49026
rect 17218 48974 17230 49026
rect 18946 48974 18958 49026
rect 19010 48974 19022 49026
rect 21298 48974 21310 49026
rect 21362 48974 21374 49026
rect 16606 48962 16658 48974
rect 21646 48962 21698 48974
rect 21870 49026 21922 49038
rect 25454 49026 25506 49038
rect 33406 49026 33458 49038
rect 23762 48974 23774 49026
rect 23826 48974 23838 49026
rect 26226 48974 26238 49026
rect 26290 48974 26302 49026
rect 27346 48974 27358 49026
rect 27410 48974 27422 49026
rect 30034 48974 30046 49026
rect 30098 48974 30110 49026
rect 30818 48974 30830 49026
rect 30882 48974 30894 49026
rect 31266 48974 31278 49026
rect 31330 48974 31342 49026
rect 33170 48974 33182 49026
rect 33234 48974 33246 49026
rect 21870 48962 21922 48974
rect 25454 48962 25506 48974
rect 33406 48962 33458 48974
rect 33630 49026 33682 49038
rect 33630 48962 33682 48974
rect 34078 49026 34130 49038
rect 35422 49026 35474 49038
rect 42814 49026 42866 49038
rect 34514 48974 34526 49026
rect 34578 48974 34590 49026
rect 34962 48974 34974 49026
rect 35026 48974 35038 49026
rect 35746 48974 35758 49026
rect 35810 48974 35822 49026
rect 39442 48974 39454 49026
rect 39506 48974 39518 49026
rect 42242 48974 42254 49026
rect 42306 48974 42318 49026
rect 34078 48962 34130 48974
rect 35422 48962 35474 48974
rect 42814 48962 42866 48974
rect 43262 49026 43314 49038
rect 43262 48962 43314 48974
rect 45950 49026 46002 49038
rect 45950 48962 46002 48974
rect 46174 49026 46226 49038
rect 46498 48974 46510 49026
rect 46562 48974 46574 49026
rect 49858 48974 49870 49026
rect 49922 48974 49934 49026
rect 46174 48962 46226 48974
rect 26462 48914 26514 48926
rect 22530 48862 22542 48914
rect 22594 48862 22606 48914
rect 22866 48862 22878 48914
rect 22930 48862 22942 48914
rect 23538 48862 23550 48914
rect 23602 48862 23614 48914
rect 26462 48850 26514 48862
rect 30270 48914 30322 48926
rect 30270 48850 30322 48862
rect 42926 48914 42978 48926
rect 42926 48850 42978 48862
rect 43934 48914 43986 48926
rect 43934 48850 43986 48862
rect 47518 48914 47570 48926
rect 47518 48850 47570 48862
rect 47742 48914 47794 48926
rect 47742 48850 47794 48862
rect 49086 48914 49138 48926
rect 49086 48850 49138 48862
rect 50878 48914 50930 48926
rect 50878 48850 50930 48862
rect 14030 48802 14082 48814
rect 14030 48738 14082 48750
rect 22206 48802 22258 48814
rect 22206 48738 22258 48750
rect 23214 48802 23266 48814
rect 23214 48738 23266 48750
rect 27134 48802 27186 48814
rect 27134 48738 27186 48750
rect 28030 48802 28082 48814
rect 28030 48738 28082 48750
rect 28590 48802 28642 48814
rect 28590 48738 28642 48750
rect 29710 48802 29762 48814
rect 29710 48738 29762 48750
rect 31390 48802 31442 48814
rect 31390 48738 31442 48750
rect 33294 48802 33346 48814
rect 33294 48738 33346 48750
rect 37774 48802 37826 48814
rect 37774 48738 37826 48750
rect 43486 48802 43538 48814
rect 43486 48738 43538 48750
rect 44158 48802 44210 48814
rect 44158 48738 44210 48750
rect 46062 48802 46114 48814
rect 46062 48738 46114 48750
rect 50990 48802 51042 48814
rect 50990 48738 51042 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 23326 48466 23378 48478
rect 21634 48414 21646 48466
rect 21698 48414 21710 48466
rect 23326 48402 23378 48414
rect 25790 48466 25842 48478
rect 34190 48466 34242 48478
rect 32162 48414 32174 48466
rect 32226 48414 32238 48466
rect 25790 48402 25842 48414
rect 34190 48402 34242 48414
rect 35646 48466 35698 48478
rect 35646 48402 35698 48414
rect 35870 48466 35922 48478
rect 35870 48402 35922 48414
rect 38446 48466 38498 48478
rect 38446 48402 38498 48414
rect 39678 48466 39730 48478
rect 39678 48402 39730 48414
rect 42366 48466 42418 48478
rect 44930 48414 44942 48466
rect 44994 48414 45006 48466
rect 42366 48402 42418 48414
rect 25902 48354 25954 48366
rect 29934 48354 29986 48366
rect 20178 48302 20190 48354
rect 20242 48302 20254 48354
rect 22642 48302 22654 48354
rect 22706 48302 22718 48354
rect 27234 48302 27246 48354
rect 27298 48302 27310 48354
rect 25902 48290 25954 48302
rect 29934 48290 29986 48302
rect 30158 48354 30210 48366
rect 34078 48354 34130 48366
rect 30482 48302 30494 48354
rect 30546 48302 30558 48354
rect 31266 48302 31278 48354
rect 31330 48302 31342 48354
rect 30158 48290 30210 48302
rect 34078 48290 34130 48302
rect 35534 48354 35586 48366
rect 37998 48354 38050 48366
rect 36418 48302 36430 48354
rect 36482 48302 36494 48354
rect 35534 48290 35586 48302
rect 37998 48290 38050 48302
rect 38558 48354 38610 48366
rect 42142 48354 42194 48366
rect 40002 48302 40014 48354
rect 40066 48302 40078 48354
rect 38558 48290 38610 48302
rect 42142 48290 42194 48302
rect 42478 48354 42530 48366
rect 45614 48354 45666 48366
rect 44034 48302 44046 48354
rect 44098 48302 44110 48354
rect 42478 48290 42530 48302
rect 45614 48290 45666 48302
rect 11230 48242 11282 48254
rect 13806 48242 13858 48254
rect 11666 48190 11678 48242
rect 11730 48190 11742 48242
rect 13346 48190 13358 48242
rect 13410 48190 13422 48242
rect 11230 48178 11282 48190
rect 13806 48178 13858 48190
rect 14142 48242 14194 48254
rect 30830 48242 30882 48254
rect 38334 48242 38386 48254
rect 15362 48190 15374 48242
rect 15426 48190 15438 48242
rect 20402 48190 20414 48242
rect 20466 48190 20478 48242
rect 21522 48190 21534 48242
rect 21586 48190 21598 48242
rect 26450 48190 26462 48242
rect 26514 48190 26526 48242
rect 27458 48190 27470 48242
rect 27522 48190 27534 48242
rect 28130 48190 28142 48242
rect 28194 48190 28206 48242
rect 28914 48190 28926 48242
rect 28978 48190 28990 48242
rect 29474 48190 29486 48242
rect 29538 48190 29550 48242
rect 31154 48190 31166 48242
rect 31218 48190 31230 48242
rect 32050 48190 32062 48242
rect 32114 48190 32126 48242
rect 36306 48190 36318 48242
rect 36370 48190 36382 48242
rect 36530 48190 36542 48242
rect 36594 48190 36606 48242
rect 37202 48190 37214 48242
rect 37266 48190 37278 48242
rect 14142 48178 14194 48190
rect 30830 48178 30882 48190
rect 38334 48178 38386 48190
rect 38894 48242 38946 48254
rect 42590 48242 42642 48254
rect 49758 48242 49810 48254
rect 39106 48190 39118 48242
rect 39170 48190 39182 48242
rect 39442 48190 39454 48242
rect 39506 48190 39518 48242
rect 40226 48190 40238 48242
rect 40290 48190 40302 48242
rect 43922 48190 43934 48242
rect 43986 48190 43998 48242
rect 44930 48190 44942 48242
rect 44994 48190 45006 48242
rect 49970 48190 49982 48242
rect 50034 48190 50046 48242
rect 38894 48178 38946 48190
rect 42590 48178 42642 48190
rect 49758 48178 49810 48190
rect 16270 48130 16322 48142
rect 15474 48078 15486 48130
rect 15538 48078 15550 48130
rect 16270 48066 16322 48078
rect 18510 48130 18562 48142
rect 18510 48066 18562 48078
rect 19294 48130 19346 48142
rect 19294 48066 19346 48078
rect 24110 48130 24162 48142
rect 24110 48066 24162 48078
rect 24782 48130 24834 48142
rect 24782 48066 24834 48078
rect 25342 48130 25394 48142
rect 25342 48066 25394 48078
rect 26910 48130 26962 48142
rect 26910 48066 26962 48078
rect 41022 48130 41074 48142
rect 50654 48130 50706 48142
rect 45714 48078 45726 48130
rect 45778 48078 45790 48130
rect 41022 48066 41074 48078
rect 50654 48066 50706 48078
rect 23214 48018 23266 48030
rect 23214 47954 23266 47966
rect 23550 48018 23602 48030
rect 23550 47954 23602 47966
rect 25678 48018 25730 48030
rect 29822 48018 29874 48030
rect 28914 47966 28926 48018
rect 28978 47966 28990 48018
rect 25678 47954 25730 47966
rect 29822 47954 29874 47966
rect 34302 48018 34354 48030
rect 34302 47954 34354 47966
rect 39342 48018 39394 48030
rect 39342 47954 39394 47966
rect 45390 48018 45442 48030
rect 45390 47954 45442 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 39790 47682 39842 47694
rect 16594 47630 16606 47682
rect 16658 47630 16670 47682
rect 25330 47630 25342 47682
rect 25394 47679 25406 47682
rect 26786 47679 26798 47682
rect 25394 47633 26798 47679
rect 25394 47630 25406 47633
rect 26786 47630 26798 47633
rect 26850 47630 26862 47682
rect 30146 47630 30158 47682
rect 30210 47630 30222 47682
rect 30930 47630 30942 47682
rect 30994 47679 31006 47682
rect 30994 47633 31439 47679
rect 30994 47630 31006 47633
rect 17614 47570 17666 47582
rect 13906 47518 13918 47570
rect 13970 47518 13982 47570
rect 16706 47518 16718 47570
rect 16770 47518 16782 47570
rect 17614 47506 17666 47518
rect 19630 47570 19682 47582
rect 19630 47506 19682 47518
rect 22318 47570 22370 47582
rect 22318 47506 22370 47518
rect 22990 47570 23042 47582
rect 22990 47506 23042 47518
rect 24334 47570 24386 47582
rect 24334 47506 24386 47518
rect 27358 47570 27410 47582
rect 31393 47570 31439 47633
rect 31602 47630 31614 47682
rect 31666 47630 31678 47682
rect 39790 47618 39842 47630
rect 49310 47570 49362 47582
rect 57934 47570 57986 47582
rect 29922 47518 29934 47570
rect 29986 47518 29998 47570
rect 31378 47518 31390 47570
rect 31442 47518 31454 47570
rect 31938 47518 31950 47570
rect 32002 47518 32014 47570
rect 37426 47518 37438 47570
rect 37490 47518 37502 47570
rect 50418 47518 50430 47570
rect 50482 47518 50494 47570
rect 27358 47506 27410 47518
rect 49310 47506 49362 47518
rect 57934 47506 57986 47518
rect 19070 47458 19122 47470
rect 13570 47406 13582 47458
rect 13634 47406 13646 47458
rect 16258 47406 16270 47458
rect 16322 47406 16334 47458
rect 17266 47406 17278 47458
rect 17330 47406 17342 47458
rect 18722 47406 18734 47458
rect 18786 47406 18798 47458
rect 19070 47394 19122 47406
rect 21534 47458 21586 47470
rect 21534 47394 21586 47406
rect 23998 47458 24050 47470
rect 23998 47394 24050 47406
rect 24446 47458 24498 47470
rect 24446 47394 24498 47406
rect 24782 47458 24834 47470
rect 27470 47458 27522 47470
rect 27010 47406 27022 47458
rect 27074 47406 27086 47458
rect 24782 47394 24834 47406
rect 27470 47394 27522 47406
rect 27582 47458 27634 47470
rect 27582 47394 27634 47406
rect 28142 47458 28194 47470
rect 36542 47458 36594 47470
rect 49534 47458 49586 47470
rect 29250 47406 29262 47458
rect 29314 47406 29326 47458
rect 30258 47406 30270 47458
rect 30322 47406 30334 47458
rect 32050 47406 32062 47458
rect 32114 47406 32126 47458
rect 37202 47406 37214 47458
rect 37266 47406 37278 47458
rect 39554 47406 39566 47458
rect 39618 47406 39630 47458
rect 39890 47406 39902 47458
rect 39954 47406 39966 47458
rect 46610 47406 46622 47458
rect 46674 47406 46686 47458
rect 50642 47406 50654 47458
rect 50706 47406 50718 47458
rect 55570 47406 55582 47458
rect 55634 47406 55646 47458
rect 28142 47394 28194 47406
rect 36542 47394 36594 47406
rect 49534 47394 49586 47406
rect 19742 47346 19794 47358
rect 18498 47294 18510 47346
rect 18562 47294 18574 47346
rect 19742 47282 19794 47294
rect 20526 47346 20578 47358
rect 20526 47282 20578 47294
rect 20638 47346 20690 47358
rect 20638 47282 20690 47294
rect 23550 47346 23602 47358
rect 23550 47282 23602 47294
rect 24222 47346 24274 47358
rect 24222 47282 24274 47294
rect 27246 47346 27298 47358
rect 27246 47282 27298 47294
rect 28254 47346 28306 47358
rect 28254 47282 28306 47294
rect 36206 47346 36258 47358
rect 36206 47282 36258 47294
rect 38110 47346 38162 47358
rect 38110 47282 38162 47294
rect 39342 47346 39394 47358
rect 39342 47282 39394 47294
rect 45502 47346 45554 47358
rect 45502 47282 45554 47294
rect 46958 47346 47010 47358
rect 46958 47282 47010 47294
rect 51326 47346 51378 47358
rect 51326 47282 51378 47294
rect 12350 47234 12402 47246
rect 12350 47170 12402 47182
rect 13022 47234 13074 47246
rect 13022 47170 13074 47182
rect 14702 47234 14754 47246
rect 14702 47170 14754 47182
rect 15598 47234 15650 47246
rect 15598 47170 15650 47182
rect 18174 47234 18226 47246
rect 18174 47170 18226 47182
rect 19518 47234 19570 47246
rect 19518 47170 19570 47182
rect 20302 47234 20354 47246
rect 20302 47170 20354 47182
rect 22766 47234 22818 47246
rect 22766 47170 22818 47182
rect 22878 47234 22930 47246
rect 22878 47170 22930 47182
rect 23326 47234 23378 47246
rect 23326 47170 23378 47182
rect 23438 47234 23490 47246
rect 23438 47170 23490 47182
rect 25342 47234 25394 47246
rect 25342 47170 25394 47182
rect 25678 47234 25730 47246
rect 25678 47170 25730 47182
rect 26126 47234 26178 47246
rect 26126 47170 26178 47182
rect 26686 47234 26738 47246
rect 26686 47170 26738 47182
rect 28030 47234 28082 47246
rect 28030 47170 28082 47182
rect 28478 47234 28530 47246
rect 28478 47170 28530 47182
rect 31166 47234 31218 47246
rect 31166 47170 31218 47182
rect 36318 47234 36370 47246
rect 36318 47170 36370 47182
rect 40126 47234 40178 47246
rect 40126 47170 40178 47182
rect 45614 47234 45666 47246
rect 45614 47170 45666 47182
rect 46846 47234 46898 47246
rect 49858 47182 49870 47234
rect 49922 47182 49934 47234
rect 46846 47170 46898 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 16046 46898 16098 46910
rect 19070 46898 19122 46910
rect 16818 46846 16830 46898
rect 16882 46846 16894 46898
rect 16046 46834 16098 46846
rect 19070 46834 19122 46846
rect 23774 46898 23826 46910
rect 23774 46834 23826 46846
rect 24222 46898 24274 46910
rect 24222 46834 24274 46846
rect 25342 46898 25394 46910
rect 25342 46834 25394 46846
rect 31278 46898 31330 46910
rect 31278 46834 31330 46846
rect 31390 46898 31442 46910
rect 31390 46834 31442 46846
rect 35422 46898 35474 46910
rect 41010 46846 41022 46898
rect 41074 46846 41086 46898
rect 35422 46834 35474 46846
rect 18062 46786 18114 46798
rect 14018 46734 14030 46786
rect 14082 46734 14094 46786
rect 14354 46734 14366 46786
rect 14418 46734 14430 46786
rect 15026 46734 15038 46786
rect 15090 46734 15102 46786
rect 18062 46722 18114 46734
rect 18846 46786 18898 46798
rect 21310 46786 21362 46798
rect 20962 46734 20974 46786
rect 21026 46734 21038 46786
rect 18846 46722 18898 46734
rect 21310 46722 21362 46734
rect 21422 46786 21474 46798
rect 23662 46786 23714 46798
rect 23090 46734 23102 46786
rect 23154 46734 23166 46786
rect 21422 46722 21474 46734
rect 23662 46722 23714 46734
rect 23886 46786 23938 46798
rect 23886 46722 23938 46734
rect 24446 46786 24498 46798
rect 24446 46722 24498 46734
rect 24558 46786 24610 46798
rect 42030 46786 42082 46798
rect 44158 46786 44210 46798
rect 35074 46734 35086 46786
rect 35138 46734 35150 46786
rect 42914 46734 42926 46786
rect 42978 46734 42990 46786
rect 24558 46722 24610 46734
rect 42030 46722 42082 46734
rect 44158 46722 44210 46734
rect 45166 46786 45218 46798
rect 51102 46786 51154 46798
rect 46498 46734 46510 46786
rect 46562 46734 46574 46786
rect 52434 46734 52446 46786
rect 52498 46734 52510 46786
rect 45166 46722 45218 46734
rect 51102 46722 51154 46734
rect 14702 46674 14754 46686
rect 17838 46674 17890 46686
rect 11666 46622 11678 46674
rect 11730 46622 11742 46674
rect 13010 46622 13022 46674
rect 13074 46622 13086 46674
rect 13794 46622 13806 46674
rect 13858 46622 13870 46674
rect 17714 46622 17726 46674
rect 17778 46622 17790 46674
rect 14702 46610 14754 46622
rect 17838 46610 17890 46622
rect 19406 46674 19458 46686
rect 21646 46674 21698 46686
rect 27246 46674 27298 46686
rect 19842 46622 19854 46674
rect 19906 46622 19918 46674
rect 20626 46622 20638 46674
rect 20690 46622 20702 46674
rect 21858 46622 21870 46674
rect 21922 46622 21934 46674
rect 22530 46622 22542 46674
rect 22594 46622 22606 46674
rect 19406 46610 19458 46622
rect 21646 46610 21698 46622
rect 27246 46610 27298 46622
rect 27694 46674 27746 46686
rect 31166 46674 31218 46686
rect 30818 46622 30830 46674
rect 30882 46622 30894 46674
rect 27694 46610 27746 46622
rect 31166 46610 31218 46622
rect 41358 46674 41410 46686
rect 41358 46610 41410 46622
rect 41806 46674 41858 46686
rect 45054 46674 45106 46686
rect 42578 46622 42590 46674
rect 42642 46622 42654 46674
rect 43138 46622 43150 46674
rect 43202 46622 43214 46674
rect 43922 46622 43934 46674
rect 43986 46622 43998 46674
rect 41806 46610 41858 46622
rect 45054 46610 45106 46622
rect 45390 46674 45442 46686
rect 50654 46674 50706 46686
rect 47506 46622 47518 46674
rect 47570 46622 47582 46674
rect 45390 46610 45442 46622
rect 50654 46610 50706 46622
rect 51326 46674 51378 46686
rect 51326 46610 51378 46622
rect 51438 46674 51490 46686
rect 51438 46610 51490 46622
rect 52894 46674 52946 46686
rect 53330 46622 53342 46674
rect 53394 46622 53406 46674
rect 52894 46610 52946 46622
rect 11230 46562 11282 46574
rect 11230 46498 11282 46510
rect 12350 46562 12402 46574
rect 12350 46498 12402 46510
rect 15486 46562 15538 46574
rect 15486 46498 15538 46510
rect 16270 46562 16322 46574
rect 16270 46498 16322 46510
rect 17950 46562 18002 46574
rect 26686 46562 26738 46574
rect 20290 46510 20302 46562
rect 20354 46510 20366 46562
rect 22642 46510 22654 46562
rect 22706 46510 22718 46562
rect 25778 46510 25790 46562
rect 25842 46510 25854 46562
rect 17950 46498 18002 46510
rect 26686 46498 26738 46510
rect 28142 46562 28194 46574
rect 28142 46498 28194 46510
rect 28702 46562 28754 46574
rect 28702 46498 28754 46510
rect 29038 46562 29090 46574
rect 29038 46498 29090 46510
rect 30494 46562 30546 46574
rect 48190 46562 48242 46574
rect 42130 46510 42142 46562
rect 42194 46510 42206 46562
rect 44594 46510 44606 46562
rect 44658 46510 44670 46562
rect 46050 46510 46062 46562
rect 46114 46510 46126 46562
rect 53106 46510 53118 46562
rect 53170 46510 53182 46562
rect 30494 46498 30546 46510
rect 48190 46498 48242 46510
rect 12686 46450 12738 46462
rect 12686 46386 12738 46398
rect 13022 46450 13074 46462
rect 13022 46386 13074 46398
rect 16494 46450 16546 46462
rect 16494 46386 16546 46398
rect 17390 46450 17442 46462
rect 17390 46386 17442 46398
rect 19182 46450 19234 46462
rect 27010 46398 27022 46450
rect 27074 46398 27086 46450
rect 19182 46386 19234 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 13694 46114 13746 46126
rect 13694 46050 13746 46062
rect 18622 46114 18674 46126
rect 18622 46050 18674 46062
rect 19966 46114 20018 46126
rect 51662 46114 51714 46126
rect 32722 46062 32734 46114
rect 32786 46062 32798 46114
rect 35858 46062 35870 46114
rect 35922 46062 35934 46114
rect 19966 46050 20018 46062
rect 51662 46050 51714 46062
rect 18286 46002 18338 46014
rect 11890 45950 11902 46002
rect 11954 45950 11966 46002
rect 12450 45950 12462 46002
rect 12514 45950 12526 46002
rect 16034 45950 16046 46002
rect 16098 45950 16110 46002
rect 35186 45950 35198 46002
rect 35250 45950 35262 46002
rect 18286 45938 18338 45950
rect 13470 45890 13522 45902
rect 14142 45890 14194 45902
rect 11554 45838 11566 45890
rect 11618 45838 11630 45890
rect 14018 45838 14030 45890
rect 14082 45838 14094 45890
rect 13470 45826 13522 45838
rect 14142 45826 14194 45838
rect 14254 45890 14306 45902
rect 14254 45826 14306 45838
rect 14366 45890 14418 45902
rect 16606 45890 16658 45902
rect 14914 45838 14926 45890
rect 14978 45838 14990 45890
rect 15474 45838 15486 45890
rect 15538 45838 15550 45890
rect 16258 45838 16270 45890
rect 16322 45838 16334 45890
rect 14366 45826 14418 45838
rect 16606 45826 16658 45838
rect 16942 45890 16994 45902
rect 16942 45826 16994 45838
rect 17390 45890 17442 45902
rect 17390 45826 17442 45838
rect 17502 45890 17554 45902
rect 17502 45826 17554 45838
rect 17614 45890 17666 45902
rect 17614 45826 17666 45838
rect 17726 45890 17778 45902
rect 19742 45890 19794 45902
rect 27022 45890 27074 45902
rect 17938 45838 17950 45890
rect 18002 45838 18014 45890
rect 20066 45838 20078 45890
rect 20130 45838 20142 45890
rect 21858 45838 21870 45890
rect 21922 45838 21934 45890
rect 23090 45838 23102 45890
rect 23154 45838 23166 45890
rect 23426 45838 23438 45890
rect 23490 45838 23502 45890
rect 23762 45838 23774 45890
rect 23826 45838 23838 45890
rect 26674 45838 26686 45890
rect 26738 45838 26750 45890
rect 17726 45826 17778 45838
rect 19742 45826 19794 45838
rect 27022 45826 27074 45838
rect 27470 45890 27522 45902
rect 27470 45826 27522 45838
rect 28366 45890 28418 45902
rect 39118 45890 39170 45902
rect 31154 45838 31166 45890
rect 31218 45838 31230 45890
rect 31602 45838 31614 45890
rect 31666 45838 31678 45890
rect 32498 45838 32510 45890
rect 32562 45838 32574 45890
rect 32834 45838 32846 45890
rect 32898 45838 32910 45890
rect 33506 45838 33518 45890
rect 33570 45838 33582 45890
rect 35074 45838 35086 45890
rect 35138 45838 35150 45890
rect 28366 45826 28418 45838
rect 39118 45826 39170 45838
rect 43822 45890 43874 45902
rect 43822 45826 43874 45838
rect 44046 45890 44098 45902
rect 44046 45826 44098 45838
rect 45390 45890 45442 45902
rect 45390 45826 45442 45838
rect 45726 45890 45778 45902
rect 45726 45826 45778 45838
rect 46510 45890 46562 45902
rect 46510 45826 46562 45838
rect 46846 45890 46898 45902
rect 46846 45826 46898 45838
rect 47070 45890 47122 45902
rect 47070 45826 47122 45838
rect 49534 45890 49586 45902
rect 50318 45890 50370 45902
rect 49858 45838 49870 45890
rect 49922 45838 49934 45890
rect 51650 45838 51662 45890
rect 51714 45838 51726 45890
rect 52882 45838 52894 45890
rect 52946 45838 52958 45890
rect 49534 45826 49586 45838
rect 50318 45826 50370 45838
rect 16718 45778 16770 45790
rect 16718 45714 16770 45726
rect 18510 45778 18562 45790
rect 27694 45778 27746 45790
rect 25218 45726 25230 45778
rect 25282 45726 25294 45778
rect 18510 45714 18562 45726
rect 27694 45714 27746 45726
rect 27806 45778 27858 45790
rect 27806 45714 27858 45726
rect 28030 45778 28082 45790
rect 28030 45714 28082 45726
rect 29262 45778 29314 45790
rect 29262 45714 29314 45726
rect 30046 45778 30098 45790
rect 31838 45778 31890 45790
rect 39454 45778 39506 45790
rect 30930 45726 30942 45778
rect 30994 45726 31006 45778
rect 33730 45726 33742 45778
rect 33794 45726 33806 45778
rect 34290 45726 34302 45778
rect 34354 45726 34366 45778
rect 38546 45726 38558 45778
rect 38610 45726 38622 45778
rect 38882 45726 38894 45778
rect 38946 45726 38958 45778
rect 30046 45714 30098 45726
rect 31838 45714 31890 45726
rect 39454 45714 39506 45726
rect 43710 45778 43762 45790
rect 43710 45714 43762 45726
rect 44270 45778 44322 45790
rect 44270 45714 44322 45726
rect 45502 45778 45554 45790
rect 45502 45714 45554 45726
rect 51326 45778 51378 45790
rect 51326 45714 51378 45726
rect 53118 45778 53170 45790
rect 53118 45714 53170 45726
rect 12910 45666 12962 45678
rect 12910 45602 12962 45614
rect 19070 45666 19122 45678
rect 19070 45602 19122 45614
rect 19518 45666 19570 45678
rect 19518 45602 19570 45614
rect 20302 45666 20354 45678
rect 20302 45602 20354 45614
rect 20750 45666 20802 45678
rect 27246 45666 27298 45678
rect 26674 45614 26686 45666
rect 26738 45614 26750 45666
rect 20750 45602 20802 45614
rect 27246 45602 27298 45614
rect 28142 45666 28194 45678
rect 28142 45602 28194 45614
rect 29710 45666 29762 45678
rect 29710 45602 29762 45614
rect 30606 45666 30658 45678
rect 40126 45666 40178 45678
rect 33954 45614 33966 45666
rect 34018 45614 34030 45666
rect 30606 45602 30658 45614
rect 40126 45602 40178 45614
rect 40462 45666 40514 45678
rect 40462 45602 40514 45614
rect 46734 45666 46786 45678
rect 46734 45602 46786 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 10558 45330 10610 45342
rect 10558 45266 10610 45278
rect 17390 45330 17442 45342
rect 17390 45266 17442 45278
rect 18398 45330 18450 45342
rect 18398 45266 18450 45278
rect 18846 45330 18898 45342
rect 18846 45266 18898 45278
rect 26462 45330 26514 45342
rect 26462 45266 26514 45278
rect 26686 45330 26738 45342
rect 26686 45266 26738 45278
rect 28030 45330 28082 45342
rect 28030 45266 28082 45278
rect 31726 45330 31778 45342
rect 31726 45266 31778 45278
rect 34638 45330 34690 45342
rect 34638 45266 34690 45278
rect 40014 45330 40066 45342
rect 40014 45266 40066 45278
rect 42702 45330 42754 45342
rect 44818 45278 44830 45330
rect 44882 45278 44894 45330
rect 42702 45266 42754 45278
rect 16718 45218 16770 45230
rect 10882 45166 10894 45218
rect 10946 45166 10958 45218
rect 16718 45154 16770 45166
rect 19966 45218 20018 45230
rect 19966 45154 20018 45166
rect 24446 45218 24498 45230
rect 29038 45218 29090 45230
rect 25330 45166 25342 45218
rect 25394 45166 25406 45218
rect 26002 45166 26014 45218
rect 26066 45166 26078 45218
rect 24446 45154 24498 45166
rect 29038 45154 29090 45166
rect 30046 45218 30098 45230
rect 37998 45218 38050 45230
rect 30818 45166 30830 45218
rect 30882 45166 30894 45218
rect 30046 45154 30098 45166
rect 37998 45154 38050 45166
rect 41918 45218 41970 45230
rect 41918 45154 41970 45166
rect 46398 45218 46450 45230
rect 46398 45154 46450 45166
rect 19854 45106 19906 45118
rect 11330 45054 11342 45106
rect 11394 45054 11406 45106
rect 11890 45054 11902 45106
rect 11954 45054 11966 45106
rect 13010 45054 13022 45106
rect 13074 45054 13086 45106
rect 14354 45054 14366 45106
rect 14418 45054 14430 45106
rect 15026 45054 15038 45106
rect 15090 45054 15102 45106
rect 16258 45054 16270 45106
rect 16322 45054 16334 45106
rect 19854 45042 19906 45054
rect 20190 45106 20242 45118
rect 24334 45106 24386 45118
rect 27022 45106 27074 45118
rect 22754 45054 22766 45106
rect 22818 45054 22830 45106
rect 23874 45054 23886 45106
rect 23938 45054 23950 45106
rect 25666 45054 25678 45106
rect 25730 45054 25742 45106
rect 20190 45042 20242 45054
rect 24334 45042 24386 45054
rect 27022 45042 27074 45054
rect 27470 45106 27522 45118
rect 34190 45106 34242 45118
rect 27794 45054 27806 45106
rect 27858 45054 27870 45106
rect 28578 45054 28590 45106
rect 28642 45054 28654 45106
rect 29474 45054 29486 45106
rect 29538 45054 29550 45106
rect 30594 45054 30606 45106
rect 30658 45054 30670 45106
rect 27470 45042 27522 45054
rect 34190 45042 34242 45054
rect 34414 45106 34466 45118
rect 34414 45042 34466 45054
rect 34862 45106 34914 45118
rect 34862 45042 34914 45054
rect 37886 45106 37938 45118
rect 37886 45042 37938 45054
rect 38222 45106 38274 45118
rect 38222 45042 38274 45054
rect 38558 45106 38610 45118
rect 39454 45106 39506 45118
rect 42254 45106 42306 45118
rect 38770 45054 38782 45106
rect 38834 45054 38846 45106
rect 39778 45054 39790 45106
rect 39842 45054 39854 45106
rect 41234 45054 41246 45106
rect 41298 45054 41310 45106
rect 38558 45042 38610 45054
rect 39454 45042 39506 45054
rect 42254 45042 42306 45054
rect 42478 45106 42530 45118
rect 46286 45106 46338 45118
rect 44594 45054 44606 45106
rect 44658 45054 44670 45106
rect 42478 45042 42530 45054
rect 46286 45042 46338 45054
rect 46622 45106 46674 45118
rect 46622 45042 46674 45054
rect 49758 45106 49810 45118
rect 49758 45042 49810 45054
rect 22094 44994 22146 45006
rect 11106 44942 11118 44994
rect 11170 44942 11182 44994
rect 14466 44942 14478 44994
rect 14530 44942 14542 44994
rect 17826 44942 17838 44994
rect 17890 44942 17902 44994
rect 22094 44930 22146 44942
rect 22654 44994 22706 45006
rect 22654 44930 22706 44942
rect 26798 44994 26850 45006
rect 26798 44930 26850 44942
rect 32286 44994 32338 45006
rect 32286 44930 32338 44942
rect 35198 44994 35250 45006
rect 42366 44994 42418 45006
rect 41010 44942 41022 44994
rect 41074 44942 41086 44994
rect 35198 44930 35250 44942
rect 42366 44930 42418 44942
rect 49534 44994 49586 45006
rect 49534 44930 49586 44942
rect 23662 44882 23714 44894
rect 23662 44818 23714 44830
rect 24446 44882 24498 44894
rect 24446 44818 24498 44830
rect 28142 44882 28194 44894
rect 31390 44882 31442 44894
rect 29698 44830 29710 44882
rect 29762 44830 29774 44882
rect 28142 44818 28194 44830
rect 31390 44818 31442 44830
rect 40126 44882 40178 44894
rect 50082 44830 50094 44882
rect 50146 44830 50158 44882
rect 40126 44818 40178 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 15822 44546 15874 44558
rect 15822 44482 15874 44494
rect 37326 44546 37378 44558
rect 37326 44482 37378 44494
rect 50878 44546 50930 44558
rect 50878 44482 50930 44494
rect 14366 44434 14418 44446
rect 12226 44382 12238 44434
rect 12290 44382 12302 44434
rect 14366 44370 14418 44382
rect 22430 44434 22482 44446
rect 22430 44370 22482 44382
rect 29262 44434 29314 44446
rect 39118 44434 39170 44446
rect 34850 44382 34862 44434
rect 34914 44382 34926 44434
rect 29262 44370 29314 44382
rect 39118 44370 39170 44382
rect 39678 44434 39730 44446
rect 57934 44434 57986 44446
rect 42690 44382 42702 44434
rect 42754 44382 42766 44434
rect 46162 44382 46174 44434
rect 46226 44382 46238 44434
rect 47506 44382 47518 44434
rect 47570 44382 47582 44434
rect 39678 44370 39730 44382
rect 57934 44370 57986 44382
rect 14590 44322 14642 44334
rect 10098 44270 10110 44322
rect 10162 44270 10174 44322
rect 10882 44270 10894 44322
rect 10946 44270 10958 44322
rect 14590 44258 14642 44270
rect 14926 44322 14978 44334
rect 14926 44258 14978 44270
rect 15150 44322 15202 44334
rect 15150 44258 15202 44270
rect 15934 44322 15986 44334
rect 21310 44322 21362 44334
rect 16930 44270 16942 44322
rect 16994 44270 17006 44322
rect 20738 44270 20750 44322
rect 20802 44270 20814 44322
rect 15934 44258 15986 44270
rect 21310 44258 21362 44270
rect 21758 44322 21810 44334
rect 35310 44322 35362 44334
rect 23650 44270 23662 44322
rect 23714 44270 23726 44322
rect 24994 44270 25006 44322
rect 25058 44270 25070 44322
rect 25330 44270 25342 44322
rect 25394 44270 25406 44322
rect 26562 44270 26574 44322
rect 26626 44270 26638 44322
rect 28242 44270 28254 44322
rect 28306 44270 28318 44322
rect 29810 44270 29822 44322
rect 29874 44270 29886 44322
rect 31154 44270 31166 44322
rect 31218 44270 31230 44322
rect 31490 44270 31502 44322
rect 31554 44270 31566 44322
rect 34626 44270 34638 44322
rect 34690 44270 34702 44322
rect 21758 44258 21810 44270
rect 35310 44258 35362 44270
rect 36990 44322 37042 44334
rect 46846 44322 46898 44334
rect 37314 44270 37326 44322
rect 37378 44270 37390 44322
rect 38658 44270 38670 44322
rect 38722 44270 38734 44322
rect 42354 44270 42366 44322
rect 42418 44270 42430 44322
rect 43474 44270 43486 44322
rect 43538 44270 43550 44322
rect 45938 44270 45950 44322
rect 46002 44270 46014 44322
rect 47394 44270 47406 44322
rect 47458 44270 47470 44322
rect 51202 44270 51214 44322
rect 51266 44270 51278 44322
rect 55570 44270 55582 44322
rect 55634 44270 55646 44322
rect 36990 44258 37042 44270
rect 46846 44258 46898 44270
rect 19630 44210 19682 44222
rect 10770 44158 10782 44210
rect 10834 44158 10846 44210
rect 17042 44158 17054 44210
rect 17106 44158 17118 44210
rect 19630 44146 19682 44158
rect 22094 44210 22146 44222
rect 39230 44210 39282 44222
rect 48302 44210 48354 44222
rect 27122 44158 27134 44210
rect 27186 44158 27198 44210
rect 31826 44158 31838 44210
rect 31890 44158 31902 44210
rect 42690 44158 42702 44210
rect 42754 44158 42766 44210
rect 22094 44146 22146 44158
rect 39230 44146 39282 44158
rect 48302 44146 48354 44158
rect 52670 44210 52722 44222
rect 52670 44146 52722 44158
rect 53006 44210 53058 44222
rect 53006 44146 53058 44158
rect 14702 44098 14754 44110
rect 10322 44046 10334 44098
rect 10386 44046 10398 44098
rect 14702 44034 14754 44046
rect 15486 44098 15538 44110
rect 15486 44034 15538 44046
rect 15710 44098 15762 44110
rect 15710 44034 15762 44046
rect 16382 44098 16434 44110
rect 16382 44034 16434 44046
rect 16494 44098 16546 44110
rect 16494 44034 16546 44046
rect 16606 44098 16658 44110
rect 22990 44098 23042 44110
rect 38334 44098 38386 44110
rect 20514 44046 20526 44098
rect 20578 44046 20590 44098
rect 26898 44046 26910 44098
rect 26962 44046 26974 44098
rect 16606 44034 16658 44046
rect 22990 44034 23042 44046
rect 38334 44034 38386 44046
rect 39006 44098 39058 44110
rect 39006 44034 39058 44046
rect 50990 44098 51042 44110
rect 50990 44034 51042 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 18846 43762 18898 43774
rect 18846 43698 18898 43710
rect 31278 43762 31330 43774
rect 31278 43698 31330 43710
rect 43038 43762 43090 43774
rect 43038 43698 43090 43710
rect 47406 43762 47458 43774
rect 47406 43698 47458 43710
rect 47630 43762 47682 43774
rect 50530 43710 50542 43762
rect 50594 43710 50606 43762
rect 47630 43698 47682 43710
rect 13582 43650 13634 43662
rect 12450 43598 12462 43650
rect 12514 43598 12526 43650
rect 13582 43586 13634 43598
rect 13694 43650 13746 43662
rect 13694 43586 13746 43598
rect 16382 43650 16434 43662
rect 16382 43586 16434 43598
rect 16830 43650 16882 43662
rect 16830 43586 16882 43598
rect 17502 43650 17554 43662
rect 17502 43586 17554 43598
rect 17614 43650 17666 43662
rect 17614 43586 17666 43598
rect 19070 43650 19122 43662
rect 19070 43586 19122 43598
rect 27246 43650 27298 43662
rect 27246 43586 27298 43598
rect 27470 43650 27522 43662
rect 27470 43586 27522 43598
rect 28590 43650 28642 43662
rect 28590 43586 28642 43598
rect 29710 43650 29762 43662
rect 29710 43586 29762 43598
rect 33854 43650 33906 43662
rect 38782 43650 38834 43662
rect 34738 43598 34750 43650
rect 34802 43598 34814 43650
rect 35746 43598 35758 43650
rect 35810 43598 35822 43650
rect 33854 43586 33906 43598
rect 38782 43586 38834 43598
rect 41022 43650 41074 43662
rect 41022 43586 41074 43598
rect 42814 43650 42866 43662
rect 42814 43586 42866 43598
rect 49758 43650 49810 43662
rect 50642 43598 50654 43650
rect 50706 43598 50718 43650
rect 49758 43586 49810 43598
rect 10222 43538 10274 43550
rect 10222 43474 10274 43486
rect 10446 43538 10498 43550
rect 10446 43474 10498 43486
rect 10894 43538 10946 43550
rect 15710 43538 15762 43550
rect 11554 43486 11566 43538
rect 11618 43486 11630 43538
rect 12114 43486 12126 43538
rect 12178 43486 12190 43538
rect 10894 43474 10946 43486
rect 15710 43474 15762 43486
rect 17726 43538 17778 43550
rect 17726 43474 17778 43486
rect 18734 43538 18786 43550
rect 18734 43474 18786 43486
rect 19518 43538 19570 43550
rect 25230 43538 25282 43550
rect 20514 43486 20526 43538
rect 20578 43486 20590 43538
rect 22194 43486 22206 43538
rect 22258 43486 22270 43538
rect 23538 43486 23550 43538
rect 23602 43486 23614 43538
rect 19518 43474 19570 43486
rect 25230 43474 25282 43486
rect 26798 43538 26850 43550
rect 26798 43474 26850 43486
rect 27582 43538 27634 43550
rect 27582 43474 27634 43486
rect 29150 43538 29202 43550
rect 29150 43474 29202 43486
rect 30270 43538 30322 43550
rect 32286 43538 32338 43550
rect 47518 43538 47570 43550
rect 30706 43486 30718 43538
rect 30770 43486 30782 43538
rect 31042 43486 31054 43538
rect 31106 43486 31118 43538
rect 34290 43486 34302 43538
rect 34354 43486 34366 43538
rect 35858 43486 35870 43538
rect 35922 43486 35934 43538
rect 38098 43486 38110 43538
rect 38162 43486 38174 43538
rect 42018 43486 42030 43538
rect 42082 43486 42094 43538
rect 44930 43486 44942 43538
rect 44994 43486 45006 43538
rect 47058 43486 47070 43538
rect 47122 43486 47134 43538
rect 50418 43486 50430 43538
rect 50482 43486 50494 43538
rect 51202 43486 51214 43538
rect 51266 43486 51278 43538
rect 52322 43486 52334 43538
rect 52386 43486 52398 43538
rect 30270 43474 30322 43486
rect 32286 43474 32338 43486
rect 47518 43474 47570 43486
rect 13022 43426 13074 43438
rect 11890 43374 11902 43426
rect 11954 43374 11966 43426
rect 13022 43362 13074 43374
rect 14590 43426 14642 43438
rect 14590 43362 14642 43374
rect 18398 43426 18450 43438
rect 18398 43362 18450 43374
rect 19294 43426 19346 43438
rect 28142 43426 28194 43438
rect 20290 43374 20302 43426
rect 20354 43374 20366 43426
rect 23874 43374 23886 43426
rect 23938 43374 23950 43426
rect 25554 43374 25566 43426
rect 25618 43374 25630 43426
rect 19294 43362 19346 43374
rect 28142 43362 28194 43374
rect 31950 43426 32002 43438
rect 39230 43426 39282 43438
rect 42366 43426 42418 43438
rect 36194 43374 36206 43426
rect 36258 43374 36270 43426
rect 37874 43374 37886 43426
rect 37938 43374 37950 43426
rect 41570 43374 41582 43426
rect 41634 43374 41646 43426
rect 31950 43362 32002 43374
rect 39230 43362 39282 43374
rect 42366 43362 42418 43374
rect 45166 43426 45218 43438
rect 45166 43362 45218 43374
rect 50990 43426 51042 43438
rect 52434 43374 52446 43426
rect 52498 43374 52510 43426
rect 50990 43362 51042 43374
rect 10894 43314 10946 43326
rect 10894 43250 10946 43262
rect 11006 43314 11058 43326
rect 11006 43250 11058 43262
rect 13694 43314 13746 43326
rect 26910 43314 26962 43326
rect 19842 43262 19854 43314
rect 19906 43262 19918 43314
rect 21746 43262 21758 43314
rect 21810 43262 21822 43314
rect 25442 43262 25454 43314
rect 25506 43262 25518 43314
rect 13694 43250 13746 43262
rect 26910 43250 26962 43262
rect 43150 43314 43202 43326
rect 43150 43250 43202 43262
rect 45278 43314 45330 43326
rect 45278 43250 45330 43262
rect 49534 43314 49586 43326
rect 49534 43250 49586 43262
rect 49870 43314 49922 43326
rect 52658 43262 52670 43314
rect 52722 43262 52734 43314
rect 49870 43250 49922 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 18846 42978 18898 42990
rect 15026 42926 15038 42978
rect 15090 42926 15102 42978
rect 17378 42926 17390 42978
rect 17442 42926 17454 42978
rect 18846 42914 18898 42926
rect 29374 42978 29426 42990
rect 29374 42914 29426 42926
rect 29710 42978 29762 42990
rect 29710 42914 29762 42926
rect 11230 42866 11282 42878
rect 16606 42866 16658 42878
rect 10098 42814 10110 42866
rect 10162 42814 10174 42866
rect 15586 42814 15598 42866
rect 15650 42814 15662 42866
rect 11230 42802 11282 42814
rect 16606 42802 16658 42814
rect 21646 42866 21698 42878
rect 23438 42866 23490 42878
rect 22530 42814 22542 42866
rect 22594 42814 22606 42866
rect 21646 42802 21698 42814
rect 23438 42802 23490 42814
rect 24558 42866 24610 42878
rect 24558 42802 24610 42814
rect 25790 42866 25842 42878
rect 25790 42802 25842 42814
rect 26574 42866 26626 42878
rect 28142 42866 28194 42878
rect 32622 42866 32674 42878
rect 27010 42814 27022 42866
rect 27074 42814 27086 42866
rect 30818 42814 30830 42866
rect 30882 42814 30894 42866
rect 31714 42814 31726 42866
rect 31778 42814 31790 42866
rect 26574 42802 26626 42814
rect 28142 42802 28194 42814
rect 32622 42802 32674 42814
rect 34302 42866 34354 42878
rect 37550 42866 37602 42878
rect 35186 42814 35198 42866
rect 35250 42814 35262 42866
rect 34302 42802 34354 42814
rect 37550 42802 37602 42814
rect 38110 42866 38162 42878
rect 43150 42866 43202 42878
rect 41794 42814 41806 42866
rect 41858 42814 41870 42866
rect 38110 42802 38162 42814
rect 43150 42802 43202 42814
rect 57934 42866 57986 42878
rect 57934 42802 57986 42814
rect 19630 42754 19682 42766
rect 10434 42702 10446 42754
rect 10498 42702 10510 42754
rect 13458 42702 13470 42754
rect 13522 42702 13534 42754
rect 15698 42702 15710 42754
rect 15762 42702 15774 42754
rect 18162 42702 18174 42754
rect 18226 42702 18238 42754
rect 18946 42702 18958 42754
rect 19010 42702 19022 42754
rect 19630 42690 19682 42702
rect 19854 42754 19906 42766
rect 19854 42690 19906 42702
rect 20302 42754 20354 42766
rect 20302 42690 20354 42702
rect 21758 42754 21810 42766
rect 21758 42690 21810 42702
rect 21982 42754 22034 42766
rect 30606 42754 30658 42766
rect 36318 42754 36370 42766
rect 24658 42702 24670 42754
rect 24722 42702 24734 42754
rect 34962 42702 34974 42754
rect 35026 42702 35038 42754
rect 21982 42690 22034 42702
rect 30606 42690 30658 42702
rect 36318 42690 36370 42702
rect 38446 42754 38498 42766
rect 38446 42690 38498 42702
rect 38558 42754 38610 42766
rect 39454 42754 39506 42766
rect 38994 42702 39006 42754
rect 39058 42702 39070 42754
rect 38558 42690 38610 42702
rect 39454 42690 39506 42702
rect 39902 42754 39954 42766
rect 39902 42690 39954 42702
rect 40014 42754 40066 42766
rect 40014 42690 40066 42702
rect 40238 42754 40290 42766
rect 45390 42754 45442 42766
rect 42018 42702 42030 42754
rect 42082 42702 42094 42754
rect 40238 42690 40290 42702
rect 45390 42690 45442 42702
rect 45502 42754 45554 42766
rect 45502 42690 45554 42702
rect 46174 42754 46226 42766
rect 46174 42690 46226 42702
rect 49198 42754 49250 42766
rect 50094 42754 50146 42766
rect 49634 42702 49646 42754
rect 49698 42702 49710 42754
rect 49198 42690 49250 42702
rect 50094 42690 50146 42702
rect 50766 42754 50818 42766
rect 50766 42690 50818 42702
rect 50878 42754 50930 42766
rect 55570 42702 55582 42754
rect 55634 42702 55646 42754
rect 50878 42690 50930 42702
rect 17166 42642 17218 42654
rect 17166 42578 17218 42590
rect 20526 42642 20578 42654
rect 20526 42578 20578 42590
rect 23662 42642 23714 42654
rect 23662 42578 23714 42590
rect 24222 42642 24274 42654
rect 24222 42578 24274 42590
rect 29150 42642 29202 42654
rect 29150 42578 29202 42590
rect 30382 42642 30434 42654
rect 30382 42578 30434 42590
rect 31390 42642 31442 42654
rect 31390 42578 31442 42590
rect 35646 42642 35698 42654
rect 35646 42578 35698 42590
rect 35982 42642 36034 42654
rect 35982 42578 36034 42590
rect 41358 42642 41410 42654
rect 41358 42578 41410 42590
rect 42702 42642 42754 42654
rect 42702 42578 42754 42590
rect 43038 42642 43090 42654
rect 43038 42578 43090 42590
rect 46734 42642 46786 42654
rect 46734 42578 46786 42590
rect 50430 42642 50482 42654
rect 50430 42578 50482 42590
rect 19742 42530 19794 42542
rect 19742 42466 19794 42478
rect 20638 42530 20690 42542
rect 20638 42466 20690 42478
rect 20862 42530 20914 42542
rect 20862 42466 20914 42478
rect 23774 42530 23826 42542
rect 23774 42466 23826 42478
rect 23998 42530 24050 42542
rect 23998 42466 24050 42478
rect 24446 42530 24498 42542
rect 24446 42466 24498 42478
rect 25230 42530 25282 42542
rect 25230 42466 25282 42478
rect 27470 42530 27522 42542
rect 27470 42466 27522 42478
rect 28590 42530 28642 42542
rect 28590 42466 28642 42478
rect 30830 42530 30882 42542
rect 30830 42466 30882 42478
rect 30942 42530 30994 42542
rect 30942 42466 30994 42478
rect 31614 42530 31666 42542
rect 31614 42466 31666 42478
rect 32174 42530 32226 42542
rect 32174 42466 32226 42478
rect 33742 42530 33794 42542
rect 33742 42466 33794 42478
rect 36094 42530 36146 42542
rect 43262 42530 43314 42542
rect 39218 42478 39230 42530
rect 39282 42478 39294 42530
rect 36094 42466 36146 42478
rect 43262 42466 43314 42478
rect 43486 42530 43538 42542
rect 43486 42466 43538 42478
rect 45614 42530 45666 42542
rect 45614 42466 45666 42478
rect 45838 42530 45890 42542
rect 45838 42466 45890 42478
rect 46510 42530 46562 42542
rect 46510 42466 46562 42478
rect 46846 42530 46898 42542
rect 46846 42466 46898 42478
rect 50654 42530 50706 42542
rect 50654 42466 50706 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 15598 42194 15650 42206
rect 15598 42130 15650 42142
rect 18286 42194 18338 42206
rect 18286 42130 18338 42142
rect 18846 42194 18898 42206
rect 26126 42194 26178 42206
rect 21634 42142 21646 42194
rect 21698 42142 21710 42194
rect 18846 42130 18898 42142
rect 26126 42130 26178 42142
rect 26350 42194 26402 42206
rect 35198 42194 35250 42206
rect 38670 42194 38722 42206
rect 27906 42142 27918 42194
rect 27970 42142 27982 42194
rect 31490 42142 31502 42194
rect 31554 42142 31566 42194
rect 35858 42142 35870 42194
rect 35922 42142 35934 42194
rect 26350 42130 26402 42142
rect 35198 42130 35250 42142
rect 38670 42130 38722 42142
rect 41470 42194 41522 42206
rect 41470 42130 41522 42142
rect 46286 42194 46338 42206
rect 47170 42142 47182 42194
rect 47234 42142 47246 42194
rect 51762 42142 51774 42194
rect 51826 42142 51838 42194
rect 46286 42130 46338 42142
rect 12014 42082 12066 42094
rect 18734 42082 18786 42094
rect 14242 42030 14254 42082
rect 14306 42030 14318 42082
rect 15810 42030 15822 42082
rect 15874 42030 15886 42082
rect 16818 42030 16830 42082
rect 16882 42030 16894 42082
rect 12014 42018 12066 42030
rect 18734 42018 18786 42030
rect 22878 42082 22930 42094
rect 34190 42082 34242 42094
rect 27346 42030 27358 42082
rect 27410 42030 27422 42082
rect 29250 42030 29262 42082
rect 29314 42030 29326 42082
rect 31714 42030 31726 42082
rect 31778 42030 31790 42082
rect 22878 42018 22930 42030
rect 34190 42018 34242 42030
rect 34414 42082 34466 42094
rect 34414 42018 34466 42030
rect 34638 42082 34690 42094
rect 34638 42018 34690 42030
rect 16046 41970 16098 41982
rect 21982 41970 22034 41982
rect 9650 41918 9662 41970
rect 9714 41918 9726 41970
rect 11554 41918 11566 41970
rect 11618 41918 11630 41970
rect 13234 41918 13246 41970
rect 13298 41918 13310 41970
rect 13906 41918 13918 41970
rect 13970 41918 13982 41970
rect 16594 41918 16606 41970
rect 16658 41918 16670 41970
rect 16046 41906 16098 41918
rect 21982 41906 22034 41918
rect 22654 41970 22706 41982
rect 22654 41906 22706 41918
rect 24222 41970 24274 41982
rect 24222 41906 24274 41918
rect 24782 41970 24834 41982
rect 24782 41906 24834 41918
rect 26014 41970 26066 41982
rect 34750 41970 34802 41982
rect 26562 41918 26574 41970
rect 26626 41918 26638 41970
rect 27010 41918 27022 41970
rect 27074 41918 27086 41970
rect 28018 41918 28030 41970
rect 28082 41918 28094 41970
rect 28690 41918 28702 41970
rect 28754 41918 28766 41970
rect 30258 41918 30270 41970
rect 30322 41918 30334 41970
rect 32162 41918 32174 41970
rect 32226 41918 32238 41970
rect 26014 41906 26066 41918
rect 34750 41906 34802 41918
rect 34862 41970 34914 41982
rect 34862 41906 34914 41918
rect 35310 41970 35362 41982
rect 35310 41906 35362 41918
rect 35534 41970 35586 41982
rect 35534 41906 35586 41918
rect 36206 41970 36258 41982
rect 45390 41970 45442 41982
rect 38994 41918 39006 41970
rect 39058 41918 39070 41970
rect 39778 41918 39790 41970
rect 39842 41918 39854 41970
rect 43810 41918 43822 41970
rect 43874 41918 43886 41970
rect 36206 41906 36258 41918
rect 45390 41906 45442 41918
rect 45614 41970 45666 41982
rect 51102 41970 51154 41982
rect 50642 41918 50654 41970
rect 50706 41918 50718 41970
rect 45614 41906 45666 41918
rect 51102 41906 51154 41918
rect 51438 41970 51490 41982
rect 51438 41906 51490 41918
rect 14030 41858 14082 41870
rect 9986 41806 9998 41858
rect 10050 41806 10062 41858
rect 14030 41794 14082 41806
rect 14814 41858 14866 41870
rect 14814 41794 14866 41806
rect 15150 41858 15202 41870
rect 19966 41858 20018 41870
rect 16146 41806 16158 41858
rect 16210 41806 16222 41858
rect 18386 41806 18398 41858
rect 18450 41806 18462 41858
rect 19842 41806 19854 41858
rect 19906 41806 19918 41858
rect 15150 41794 15202 41806
rect 15262 41746 15314 41758
rect 15262 41682 15314 41694
rect 18062 41746 18114 41758
rect 18062 41682 18114 41694
rect 18846 41746 18898 41758
rect 19857 41743 19903 41806
rect 19966 41794 20018 41806
rect 20414 41858 20466 41870
rect 20414 41794 20466 41806
rect 20974 41858 21026 41870
rect 20974 41794 21026 41806
rect 21422 41858 21474 41870
rect 25566 41858 25618 41870
rect 33182 41858 33234 41870
rect 23202 41806 23214 41858
rect 23266 41806 23278 41858
rect 26450 41806 26462 41858
rect 26514 41806 26526 41858
rect 21422 41794 21474 41806
rect 25566 41794 25618 41806
rect 33182 41794 33234 41806
rect 33630 41858 33682 41870
rect 46622 41858 46674 41870
rect 39666 41806 39678 41858
rect 39730 41806 39742 41858
rect 43922 41806 43934 41858
rect 43986 41806 43998 41858
rect 50194 41806 50206 41858
rect 50258 41806 50270 41858
rect 33630 41794 33682 41806
rect 46622 41794 46674 41806
rect 24558 41746 24610 41758
rect 45838 41746 45890 41758
rect 21298 41743 21310 41746
rect 19857 41697 21310 41743
rect 21298 41694 21310 41697
rect 21362 41694 21374 41746
rect 39890 41694 39902 41746
rect 39954 41694 39966 41746
rect 44482 41694 44494 41746
rect 44546 41694 44558 41746
rect 18846 41682 18898 41694
rect 24558 41682 24610 41694
rect 45838 41682 45890 41694
rect 46846 41746 46898 41758
rect 46846 41682 46898 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 14926 41410 14978 41422
rect 14926 41346 14978 41358
rect 18846 41410 18898 41422
rect 36206 41410 36258 41422
rect 19170 41358 19182 41410
rect 19234 41358 19246 41410
rect 18846 41346 18898 41358
rect 36206 41346 36258 41358
rect 45390 41410 45442 41422
rect 45390 41346 45442 41358
rect 1710 41298 1762 41310
rect 1710 41234 1762 41246
rect 8878 41298 8930 41310
rect 8878 41234 8930 41246
rect 9886 41298 9938 41310
rect 9886 41234 9938 41246
rect 10222 41298 10274 41310
rect 10222 41234 10274 41246
rect 11342 41298 11394 41310
rect 11342 41234 11394 41246
rect 15262 41298 15314 41310
rect 15262 41234 15314 41246
rect 16270 41298 16322 41310
rect 16270 41234 16322 41246
rect 18286 41298 18338 41310
rect 18286 41234 18338 41246
rect 21534 41298 21586 41310
rect 21534 41234 21586 41246
rect 22094 41298 22146 41310
rect 22094 41234 22146 41246
rect 24894 41298 24946 41310
rect 24894 41234 24946 41246
rect 27470 41298 27522 41310
rect 30382 41298 30434 41310
rect 44830 41298 44882 41310
rect 57934 41298 57986 41310
rect 29362 41246 29374 41298
rect 29426 41246 29438 41298
rect 32386 41246 32398 41298
rect 32450 41246 32462 41298
rect 34290 41246 34302 41298
rect 34354 41246 34366 41298
rect 35746 41246 35758 41298
rect 35810 41246 35822 41298
rect 39106 41246 39118 41298
rect 39170 41246 39182 41298
rect 45938 41246 45950 41298
rect 46002 41246 46014 41298
rect 49522 41246 49534 41298
rect 49586 41246 49598 41298
rect 27470 41234 27522 41246
rect 30382 41234 30434 41246
rect 44830 41234 44882 41246
rect 57934 41234 57986 41246
rect 10782 41186 10834 41198
rect 12350 41186 12402 41198
rect 16830 41186 16882 41198
rect 11778 41134 11790 41186
rect 11842 41134 11854 41186
rect 13458 41134 13470 41186
rect 13522 41134 13534 41186
rect 14578 41134 14590 41186
rect 14642 41134 14654 41186
rect 10782 41122 10834 41134
rect 12350 41122 12402 41134
rect 16830 41122 16882 41134
rect 18622 41186 18674 41198
rect 25006 41186 25058 41198
rect 28030 41186 28082 41198
rect 45054 41186 45106 41198
rect 22418 41134 22430 41186
rect 22482 41134 22494 41186
rect 24658 41134 24670 41186
rect 24722 41134 24734 41186
rect 26002 41134 26014 41186
rect 26066 41134 26078 41186
rect 27010 41134 27022 41186
rect 27074 41134 27086 41186
rect 28466 41134 28478 41186
rect 28530 41134 28542 41186
rect 31042 41134 31054 41186
rect 31106 41134 31118 41186
rect 32162 41134 32174 41186
rect 32226 41134 32238 41186
rect 32498 41134 32510 41186
rect 32562 41134 32574 41186
rect 33506 41134 33518 41186
rect 33570 41134 33582 41186
rect 34066 41134 34078 41186
rect 34130 41134 34142 41186
rect 35858 41134 35870 41186
rect 35922 41134 35934 41186
rect 47394 41134 47406 41186
rect 47458 41134 47470 41186
rect 48402 41134 48414 41186
rect 48466 41134 48478 41186
rect 49186 41134 49198 41186
rect 49250 41134 49262 41186
rect 55570 41134 55582 41186
rect 55634 41134 55646 41186
rect 18622 41122 18674 41134
rect 25006 41122 25058 41134
rect 28030 41122 28082 41134
rect 45054 41122 45106 41134
rect 8990 41074 9042 41086
rect 19518 41074 19570 41086
rect 12674 41022 12686 41074
rect 12738 41022 12750 41074
rect 13570 41022 13582 41074
rect 13634 41022 13646 41074
rect 8990 41010 9042 41022
rect 19518 41010 19570 41022
rect 19742 41074 19794 41086
rect 30494 41074 30546 41086
rect 35086 41074 35138 41086
rect 22306 41022 22318 41074
rect 22370 41022 22382 41074
rect 30818 41022 30830 41074
rect 30882 41022 30894 41074
rect 31490 41022 31502 41074
rect 31554 41022 31566 41074
rect 33058 41022 33070 41074
rect 33122 41022 33134 41074
rect 34402 41022 34414 41074
rect 34466 41022 34478 41074
rect 19742 41010 19794 41022
rect 30494 41010 30546 41022
rect 35086 41010 35138 41022
rect 35534 41074 35586 41086
rect 35534 41010 35586 41022
rect 36318 41074 36370 41086
rect 48078 41074 48130 41086
rect 46386 41022 46398 41074
rect 46450 41022 46462 41074
rect 49858 41022 49870 41074
rect 49922 41022 49934 41074
rect 36318 41010 36370 41022
rect 48078 41010 48130 41022
rect 8766 40962 8818 40974
rect 8766 40898 8818 40910
rect 9326 40962 9378 40974
rect 15038 40962 15090 40974
rect 12002 40910 12014 40962
rect 12066 40910 12078 40962
rect 14466 40910 14478 40962
rect 14530 40910 14542 40962
rect 9326 40898 9378 40910
rect 15038 40898 15090 40910
rect 19630 40962 19682 40974
rect 19630 40898 19682 40910
rect 20302 40962 20354 40974
rect 20302 40898 20354 40910
rect 20750 40962 20802 40974
rect 20750 40898 20802 40910
rect 29822 40962 29874 40974
rect 29822 40898 29874 40910
rect 30270 40962 30322 40974
rect 30270 40898 30322 40910
rect 39566 40962 39618 40974
rect 39566 40898 39618 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 15262 40626 15314 40638
rect 15262 40562 15314 40574
rect 15486 40626 15538 40638
rect 15486 40562 15538 40574
rect 15710 40626 15762 40638
rect 15710 40562 15762 40574
rect 16718 40626 16770 40638
rect 27246 40626 27298 40638
rect 16718 40562 16770 40574
rect 20078 40570 20130 40582
rect 26226 40574 26238 40626
rect 26290 40574 26302 40626
rect 10670 40514 10722 40526
rect 16270 40514 16322 40526
rect 11106 40462 11118 40514
rect 11170 40462 11182 40514
rect 13234 40462 13246 40514
rect 13298 40462 13310 40514
rect 14802 40462 14814 40514
rect 14866 40462 14878 40514
rect 10670 40450 10722 40462
rect 16270 40450 16322 40462
rect 16494 40514 16546 40526
rect 16494 40450 16546 40462
rect 17726 40514 17778 40526
rect 18286 40514 18338 40526
rect 27246 40562 27298 40574
rect 27470 40626 27522 40638
rect 27470 40562 27522 40574
rect 35646 40626 35698 40638
rect 35646 40562 35698 40574
rect 43486 40626 43538 40638
rect 50418 40574 50430 40626
rect 50482 40574 50494 40626
rect 43486 40562 43538 40574
rect 18050 40462 18062 40514
rect 18114 40462 18126 40514
rect 18722 40462 18734 40514
rect 18786 40462 18798 40514
rect 20078 40506 20130 40518
rect 26798 40514 26850 40526
rect 21522 40462 21534 40514
rect 21586 40462 21598 40514
rect 25330 40462 25342 40514
rect 25394 40462 25406 40514
rect 17726 40450 17778 40462
rect 18286 40450 18338 40462
rect 26798 40450 26850 40462
rect 34302 40514 34354 40526
rect 36530 40462 36542 40514
rect 36594 40462 36606 40514
rect 38994 40462 39006 40514
rect 39058 40462 39070 40514
rect 39442 40462 39454 40514
rect 39506 40462 39518 40514
rect 41234 40462 41246 40514
rect 41298 40462 41310 40514
rect 34302 40450 34354 40462
rect 16830 40402 16882 40414
rect 19854 40402 19906 40414
rect 27582 40402 27634 40414
rect 44046 40402 44098 40414
rect 49758 40402 49810 40414
rect 10210 40350 10222 40402
rect 10274 40350 10286 40402
rect 10994 40350 11006 40402
rect 11058 40350 11070 40402
rect 13346 40350 13358 40402
rect 13410 40350 13422 40402
rect 13682 40350 13694 40402
rect 13746 40350 13758 40402
rect 14242 40350 14254 40402
rect 14306 40350 14318 40402
rect 19170 40350 19182 40402
rect 19234 40350 19246 40402
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 20626 40350 20638 40402
rect 20690 40350 20702 40402
rect 21186 40350 21198 40402
rect 21250 40350 21262 40402
rect 24098 40350 24110 40402
rect 24162 40350 24174 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 25218 40350 25230 40402
rect 25282 40350 25294 40402
rect 26114 40350 26126 40402
rect 26178 40350 26190 40402
rect 27906 40350 27918 40402
rect 27970 40350 27982 40402
rect 28690 40350 28702 40402
rect 28754 40350 28766 40402
rect 29810 40350 29822 40402
rect 29874 40350 29886 40402
rect 30930 40350 30942 40402
rect 30994 40350 31006 40402
rect 32274 40350 32286 40402
rect 32338 40350 32350 40402
rect 33282 40350 33294 40402
rect 33346 40350 33358 40402
rect 37762 40350 37774 40402
rect 37826 40350 37838 40402
rect 39106 40350 39118 40402
rect 39170 40350 39182 40402
rect 41570 40350 41582 40402
rect 41634 40350 41646 40402
rect 42466 40350 42478 40402
rect 42530 40350 42542 40402
rect 49074 40350 49086 40402
rect 49138 40350 49150 40402
rect 49522 40350 49534 40402
rect 49586 40350 49598 40402
rect 16830 40338 16882 40350
rect 19854 40338 19906 40350
rect 27582 40338 27634 40350
rect 44046 40338 44098 40350
rect 49758 40338 49810 40350
rect 50094 40402 50146 40414
rect 50094 40338 50146 40350
rect 15598 40290 15650 40302
rect 14690 40238 14702 40290
rect 14754 40238 14766 40290
rect 15598 40226 15650 40238
rect 17390 40290 17442 40302
rect 17390 40226 17442 40238
rect 17502 40290 17554 40302
rect 27022 40290 27074 40302
rect 18386 40238 18398 40290
rect 18450 40238 18462 40290
rect 18946 40238 18958 40290
rect 19010 40238 19022 40290
rect 20178 40238 20190 40290
rect 20242 40238 20254 40290
rect 22418 40238 22430 40290
rect 22482 40238 22494 40290
rect 26674 40238 26686 40290
rect 26738 40238 26750 40290
rect 17502 40226 17554 40238
rect 27022 40226 27074 40238
rect 35086 40290 35138 40302
rect 38446 40290 38498 40302
rect 36306 40238 36318 40290
rect 36370 40238 36382 40290
rect 35086 40226 35138 40238
rect 38446 40226 38498 40238
rect 43150 40290 43202 40302
rect 43150 40226 43202 40238
rect 31826 40126 31838 40178
rect 31890 40126 31902 40178
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 37550 39842 37602 39854
rect 16818 39790 16830 39842
rect 16882 39790 16894 39842
rect 34178 39790 34190 39842
rect 34242 39790 34254 39842
rect 37550 39778 37602 39790
rect 45726 39842 45778 39854
rect 45726 39778 45778 39790
rect 9102 39730 9154 39742
rect 11342 39730 11394 39742
rect 9874 39678 9886 39730
rect 9938 39678 9950 39730
rect 9102 39666 9154 39678
rect 11342 39666 11394 39678
rect 12798 39730 12850 39742
rect 14478 39730 14530 39742
rect 13570 39678 13582 39730
rect 13634 39678 13646 39730
rect 12798 39666 12850 39678
rect 14478 39666 14530 39678
rect 19406 39730 19458 39742
rect 19406 39666 19458 39678
rect 19966 39730 20018 39742
rect 25342 39730 25394 39742
rect 30830 39730 30882 39742
rect 22754 39678 22766 39730
rect 22818 39678 22830 39730
rect 24098 39678 24110 39730
rect 24162 39678 24174 39730
rect 28466 39678 28478 39730
rect 28530 39678 28542 39730
rect 19966 39666 20018 39678
rect 25342 39666 25394 39678
rect 30830 39666 30882 39678
rect 38222 39730 38274 39742
rect 39554 39678 39566 39730
rect 39618 39678 39630 39730
rect 38222 39666 38274 39678
rect 8542 39618 8594 39630
rect 8542 39554 8594 39566
rect 9438 39618 9490 39630
rect 12686 39618 12738 39630
rect 11778 39566 11790 39618
rect 11842 39566 11854 39618
rect 9438 39554 9490 39566
rect 12686 39554 12738 39566
rect 12910 39618 12962 39630
rect 19182 39618 19234 39630
rect 15138 39566 15150 39618
rect 15202 39566 15214 39618
rect 16370 39566 16382 39618
rect 16434 39566 16446 39618
rect 17266 39566 17278 39618
rect 17330 39566 17342 39618
rect 18050 39566 18062 39618
rect 18114 39566 18126 39618
rect 12910 39554 12962 39566
rect 19182 39554 19234 39566
rect 20190 39618 20242 39630
rect 21646 39618 21698 39630
rect 25566 39618 25618 39630
rect 20514 39566 20526 39618
rect 20578 39566 20590 39618
rect 23874 39566 23886 39618
rect 23938 39566 23950 39618
rect 24210 39566 24222 39618
rect 24274 39566 24286 39618
rect 20190 39554 20242 39566
rect 21646 39554 21698 39566
rect 25566 39554 25618 39566
rect 25790 39618 25842 39630
rect 29262 39618 29314 39630
rect 26338 39566 26350 39618
rect 26402 39566 26414 39618
rect 27346 39566 27358 39618
rect 27410 39566 27422 39618
rect 27570 39566 27582 39618
rect 27634 39566 27646 39618
rect 28354 39566 28366 39618
rect 28418 39566 28430 39618
rect 25790 39554 25842 39566
rect 29262 39554 29314 39566
rect 29598 39618 29650 39630
rect 29598 39554 29650 39566
rect 30382 39618 30434 39630
rect 30382 39554 30434 39566
rect 31166 39618 31218 39630
rect 36318 39618 36370 39630
rect 41582 39618 41634 39630
rect 31378 39566 31390 39618
rect 31442 39566 31454 39618
rect 32946 39566 32958 39618
rect 33010 39566 33022 39618
rect 33170 39566 33182 39618
rect 33234 39566 33246 39618
rect 35970 39566 35982 39618
rect 36034 39566 36046 39618
rect 37202 39566 37214 39618
rect 37266 39566 37278 39618
rect 38546 39566 38558 39618
rect 38610 39566 38622 39618
rect 39106 39566 39118 39618
rect 39170 39566 39182 39618
rect 40562 39566 40574 39618
rect 40626 39566 40638 39618
rect 41122 39566 41134 39618
rect 41186 39566 41198 39618
rect 31166 39554 31218 39566
rect 36318 39554 36370 39566
rect 41582 39554 41634 39566
rect 42142 39618 42194 39630
rect 42142 39554 42194 39566
rect 42366 39618 42418 39630
rect 43374 39618 43426 39630
rect 43138 39566 43150 39618
rect 43202 39566 43214 39618
rect 42366 39554 42418 39566
rect 43374 39554 43426 39566
rect 43486 39618 43538 39630
rect 45390 39618 45442 39630
rect 46622 39618 46674 39630
rect 43922 39566 43934 39618
rect 43986 39566 43998 39618
rect 46386 39566 46398 39618
rect 46450 39566 46462 39618
rect 43486 39554 43538 39566
rect 45390 39554 45442 39566
rect 46622 39554 46674 39566
rect 46846 39618 46898 39630
rect 46846 39554 46898 39566
rect 18958 39506 19010 39518
rect 12002 39454 12014 39506
rect 12066 39454 12078 39506
rect 17826 39454 17838 39506
rect 17890 39454 17902 39506
rect 18958 39442 19010 39454
rect 19518 39506 19570 39518
rect 19518 39442 19570 39454
rect 20750 39506 20802 39518
rect 20750 39442 20802 39454
rect 21310 39506 21362 39518
rect 21310 39442 21362 39454
rect 21422 39506 21474 39518
rect 25230 39506 25282 39518
rect 29374 39506 29426 39518
rect 24882 39454 24894 39506
rect 24946 39454 24958 39506
rect 26114 39454 26126 39506
rect 26178 39454 26190 39506
rect 21422 39442 21474 39454
rect 25230 39442 25282 39454
rect 29374 39442 29426 39454
rect 36430 39506 36482 39518
rect 36430 39442 36482 39454
rect 37438 39506 37490 39518
rect 42702 39506 42754 39518
rect 39218 39454 39230 39506
rect 39282 39454 39294 39506
rect 40226 39454 40238 39506
rect 40290 39454 40302 39506
rect 37438 39442 37490 39454
rect 42702 39442 42754 39454
rect 45166 39506 45218 39518
rect 45166 39442 45218 39454
rect 10782 39394 10834 39406
rect 10782 39330 10834 39342
rect 12462 39394 12514 39406
rect 12462 39330 12514 39342
rect 14030 39394 14082 39406
rect 14030 39330 14082 39342
rect 20862 39394 20914 39406
rect 20862 39330 20914 39342
rect 23214 39394 23266 39406
rect 23214 39330 23266 39342
rect 26910 39394 26962 39406
rect 26910 39330 26962 39342
rect 29822 39394 29874 39406
rect 41470 39394 41522 39406
rect 41010 39342 41022 39394
rect 41074 39342 41086 39394
rect 29822 39330 29874 39342
rect 41470 39330 41522 39342
rect 41694 39394 41746 39406
rect 41694 39330 41746 39342
rect 46510 39394 46562 39406
rect 46510 39330 46562 39342
rect 58158 39394 58210 39406
rect 58158 39330 58210 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 8654 39058 8706 39070
rect 8654 38994 8706 39006
rect 11454 39058 11506 39070
rect 11454 38994 11506 39006
rect 14590 39058 14642 39070
rect 17726 39058 17778 39070
rect 17378 39006 17390 39058
rect 17442 39006 17454 39058
rect 14590 38994 14642 39006
rect 17726 38994 17778 39006
rect 22766 39058 22818 39070
rect 22766 38994 22818 39006
rect 29598 39058 29650 39070
rect 29598 38994 29650 39006
rect 31166 39058 31218 39070
rect 31166 38994 31218 39006
rect 31278 39058 31330 39070
rect 31278 38994 31330 39006
rect 33294 39058 33346 39070
rect 33294 38994 33346 39006
rect 34414 39058 34466 39070
rect 34414 38994 34466 39006
rect 39790 39058 39842 39070
rect 39790 38994 39842 39006
rect 41246 39058 41298 39070
rect 41246 38994 41298 39006
rect 41694 39058 41746 39070
rect 41694 38994 41746 39006
rect 42142 39058 42194 39070
rect 42142 38994 42194 39006
rect 46286 39058 46338 39070
rect 46286 38994 46338 39006
rect 10894 38946 10946 38958
rect 15150 38946 15202 38958
rect 20862 38946 20914 38958
rect 33518 38946 33570 38958
rect 12114 38894 12126 38946
rect 12178 38894 12190 38946
rect 16706 38894 16718 38946
rect 16770 38894 16782 38946
rect 24098 38894 24110 38946
rect 24162 38894 24174 38946
rect 29138 38894 29150 38946
rect 29202 38894 29214 38946
rect 30034 38894 30046 38946
rect 30098 38894 30110 38946
rect 10894 38882 10946 38894
rect 15150 38882 15202 38894
rect 20862 38882 20914 38894
rect 33518 38882 33570 38894
rect 42254 38946 42306 38958
rect 58158 38946 58210 38958
rect 43026 38894 43038 38946
rect 43090 38894 43102 38946
rect 47506 38894 47518 38946
rect 47570 38894 47582 38946
rect 42254 38882 42306 38894
rect 58158 38882 58210 38894
rect 19966 38834 20018 38846
rect 22990 38834 23042 38846
rect 10434 38782 10446 38834
rect 10498 38782 10510 38834
rect 11890 38782 11902 38834
rect 11954 38782 11966 38834
rect 13458 38782 13470 38834
rect 13522 38782 13534 38834
rect 15698 38782 15710 38834
rect 15762 38782 15774 38834
rect 16146 38782 16158 38834
rect 16210 38782 16222 38834
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 21410 38782 21422 38834
rect 21474 38782 21486 38834
rect 19966 38770 20018 38782
rect 22990 38770 23042 38782
rect 23438 38834 23490 38846
rect 23438 38770 23490 38782
rect 23662 38834 23714 38846
rect 31054 38834 31106 38846
rect 45838 38834 45890 38846
rect 23986 38782 23998 38834
rect 24050 38782 24062 38834
rect 26338 38782 26350 38834
rect 26402 38782 26414 38834
rect 27794 38782 27806 38834
rect 27858 38782 27870 38834
rect 28130 38782 28142 38834
rect 28194 38782 28206 38834
rect 30594 38782 30606 38834
rect 30658 38782 30670 38834
rect 31602 38782 31614 38834
rect 31666 38782 31678 38834
rect 34626 38782 34638 38834
rect 34690 38782 34702 38834
rect 43138 38782 43150 38834
rect 43202 38782 43214 38834
rect 43474 38782 43486 38834
rect 43538 38782 43550 38834
rect 23662 38770 23714 38782
rect 31054 38770 31106 38782
rect 45838 38770 45890 38782
rect 46398 38834 46450 38846
rect 46398 38770 46450 38782
rect 46510 38834 46562 38846
rect 46834 38782 46846 38834
rect 46898 38782 46910 38834
rect 47394 38782 47406 38834
rect 47458 38782 47470 38834
rect 46510 38770 46562 38782
rect 8766 38722 8818 38734
rect 23214 38722 23266 38734
rect 25342 38722 25394 38734
rect 33406 38722 33458 38734
rect 13234 38670 13246 38722
rect 13298 38670 13310 38722
rect 16034 38670 16046 38722
rect 16098 38670 16110 38722
rect 21522 38670 21534 38722
rect 21586 38670 21598 38722
rect 24658 38670 24670 38722
rect 24722 38670 24734 38722
rect 30258 38670 30270 38722
rect 30322 38670 30334 38722
rect 8766 38658 8818 38670
rect 23214 38658 23266 38670
rect 25342 38658 25394 38670
rect 33406 38658 33458 38670
rect 41582 38722 41634 38734
rect 43250 38670 43262 38722
rect 43314 38670 43326 38722
rect 47842 38670 47854 38722
rect 47906 38670 47918 38722
rect 41582 38658 41634 38670
rect 34302 38610 34354 38622
rect 34302 38546 34354 38558
rect 42142 38610 42194 38622
rect 42142 38546 42194 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 15934 38274 15986 38286
rect 15934 38210 15986 38222
rect 23886 38274 23938 38286
rect 23886 38210 23938 38222
rect 29710 38274 29762 38286
rect 29710 38210 29762 38222
rect 37550 38274 37602 38286
rect 37550 38210 37602 38222
rect 37774 38274 37826 38286
rect 37774 38210 37826 38222
rect 12910 38162 12962 38174
rect 12910 38098 12962 38110
rect 21646 38162 21698 38174
rect 21646 38098 21698 38110
rect 22878 38162 22930 38174
rect 26014 38162 26066 38174
rect 31166 38162 31218 38174
rect 46846 38162 46898 38174
rect 24994 38110 25006 38162
rect 25058 38110 25070 38162
rect 28242 38110 28254 38162
rect 28306 38110 28318 38162
rect 32274 38110 32286 38162
rect 32338 38110 32350 38162
rect 22878 38098 22930 38110
rect 26014 38098 26066 38110
rect 31166 38098 31218 38110
rect 46846 38098 46898 38110
rect 57934 38162 57986 38174
rect 57934 38098 57986 38110
rect 9662 38050 9714 38062
rect 12350 38050 12402 38062
rect 10994 37998 11006 38050
rect 11058 37998 11070 38050
rect 9662 37986 9714 37998
rect 12350 37986 12402 37998
rect 13806 38050 13858 38062
rect 13806 37986 13858 37998
rect 14030 38050 14082 38062
rect 19294 38050 19346 38062
rect 24110 38050 24162 38062
rect 25118 38050 25170 38062
rect 14466 37998 14478 38050
rect 14530 37998 14542 38050
rect 16482 37998 16494 38050
rect 16546 37998 16558 38050
rect 17154 37998 17166 38050
rect 17218 37998 17230 38050
rect 19506 37998 19518 38050
rect 19570 37998 19582 38050
rect 24882 37998 24894 38050
rect 24946 37998 24958 38050
rect 14030 37986 14082 37998
rect 19294 37986 19346 37998
rect 24110 37986 24162 37998
rect 25118 37986 25170 37998
rect 25342 38050 25394 38062
rect 31614 38050 31666 38062
rect 32846 38050 32898 38062
rect 26114 37998 26126 38050
rect 26178 37998 26190 38050
rect 27906 37998 27918 38050
rect 27970 37998 27982 38050
rect 29586 37998 29598 38050
rect 29650 37998 29662 38050
rect 32610 37998 32622 38050
rect 32674 37998 32686 38050
rect 25342 37986 25394 37998
rect 31614 37986 31666 37998
rect 32846 37986 32898 37998
rect 33182 38050 33234 38062
rect 33182 37986 33234 37998
rect 33406 38050 33458 38062
rect 34526 38050 34578 38062
rect 33954 37998 33966 38050
rect 34018 37998 34030 38050
rect 33406 37986 33458 37998
rect 34526 37986 34578 37998
rect 35086 38050 35138 38062
rect 35086 37986 35138 37998
rect 35198 38050 35250 38062
rect 35198 37986 35250 37998
rect 35422 38050 35474 38062
rect 35422 37986 35474 37998
rect 42814 38050 42866 38062
rect 48178 37998 48190 38050
rect 48242 37998 48254 38050
rect 55570 37998 55582 38050
rect 55634 37998 55646 38050
rect 42814 37986 42866 37998
rect 12126 37938 12178 37950
rect 19630 37938 19682 37950
rect 11106 37886 11118 37938
rect 11170 37886 11182 37938
rect 11442 37886 11454 37938
rect 11506 37886 11518 37938
rect 16594 37886 16606 37938
rect 16658 37886 16670 37938
rect 17378 37886 17390 37938
rect 17442 37886 17454 37938
rect 12126 37874 12178 37886
rect 19630 37874 19682 37886
rect 24334 37938 24386 37950
rect 24334 37874 24386 37886
rect 25566 37938 25618 37950
rect 25566 37874 25618 37886
rect 25902 37938 25954 37950
rect 25902 37874 25954 37886
rect 29262 37938 29314 37950
rect 31950 37938 32002 37950
rect 29698 37886 29710 37938
rect 29762 37886 29774 37938
rect 29262 37874 29314 37886
rect 31950 37874 32002 37886
rect 34638 37938 34690 37950
rect 34638 37874 34690 37886
rect 34974 37938 35026 37950
rect 34974 37874 35026 37886
rect 36990 37938 37042 37950
rect 36990 37874 37042 37886
rect 37886 37938 37938 37950
rect 37886 37874 37938 37886
rect 42478 37938 42530 37950
rect 48862 37938 48914 37950
rect 47170 37886 47182 37938
rect 47234 37886 47246 37938
rect 42478 37874 42530 37886
rect 48862 37874 48914 37886
rect 49198 37938 49250 37950
rect 49198 37874 49250 37886
rect 49534 37938 49586 37950
rect 49534 37874 49586 37886
rect 1710 37826 1762 37838
rect 1710 37762 1762 37774
rect 9102 37826 9154 37838
rect 9102 37762 9154 37774
rect 22206 37826 22258 37838
rect 22206 37762 22258 37774
rect 23214 37826 23266 37838
rect 23214 37762 23266 37774
rect 23550 37826 23602 37838
rect 23550 37762 23602 37774
rect 23774 37826 23826 37838
rect 23774 37762 23826 37774
rect 24446 37826 24498 37838
rect 24446 37762 24498 37774
rect 24670 37826 24722 37838
rect 24670 37762 24722 37774
rect 26350 37826 26402 37838
rect 26350 37762 26402 37774
rect 26798 37826 26850 37838
rect 26798 37762 26850 37774
rect 27470 37826 27522 37838
rect 27470 37762 27522 37774
rect 30718 37826 30770 37838
rect 30718 37762 30770 37774
rect 31726 37826 31778 37838
rect 31726 37762 31778 37774
rect 37214 37826 37266 37838
rect 37214 37762 37266 37774
rect 37438 37826 37490 37838
rect 37438 37762 37490 37774
rect 42590 37826 42642 37838
rect 42590 37762 42642 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 20414 37490 20466 37502
rect 18050 37438 18062 37490
rect 18114 37438 18126 37490
rect 20414 37426 20466 37438
rect 34302 37490 34354 37502
rect 34302 37426 34354 37438
rect 35646 37490 35698 37502
rect 35646 37426 35698 37438
rect 37214 37490 37266 37502
rect 43934 37490 43986 37502
rect 41906 37438 41918 37490
rect 41970 37438 41982 37490
rect 47282 37438 47294 37490
rect 47346 37438 47358 37490
rect 37214 37426 37266 37438
rect 43934 37426 43986 37438
rect 18958 37378 19010 37390
rect 36878 37378 36930 37390
rect 8978 37326 8990 37378
rect 9042 37326 9054 37378
rect 12450 37326 12462 37378
rect 12514 37326 12526 37378
rect 21186 37326 21198 37378
rect 21250 37326 21262 37378
rect 25554 37326 25566 37378
rect 25618 37326 25630 37378
rect 18958 37314 19010 37326
rect 36878 37314 36930 37326
rect 36990 37378 37042 37390
rect 36990 37314 37042 37326
rect 38558 37378 38610 37390
rect 38558 37314 38610 37326
rect 39342 37378 39394 37390
rect 46734 37378 46786 37390
rect 41122 37326 41134 37378
rect 41186 37326 41198 37378
rect 39342 37314 39394 37326
rect 46734 37314 46786 37326
rect 18174 37266 18226 37278
rect 7858 37214 7870 37266
rect 7922 37214 7934 37266
rect 8306 37214 8318 37266
rect 8370 37214 8382 37266
rect 9650 37214 9662 37266
rect 9714 37214 9726 37266
rect 10882 37214 10894 37266
rect 10946 37214 10958 37266
rect 12786 37214 12798 37266
rect 12850 37214 12862 37266
rect 13794 37214 13806 37266
rect 13858 37214 13870 37266
rect 16034 37214 16046 37266
rect 16098 37214 16110 37266
rect 18174 37202 18226 37214
rect 19854 37266 19906 37278
rect 29262 37266 29314 37278
rect 31278 37266 31330 37278
rect 21858 37214 21870 37266
rect 21922 37214 21934 37266
rect 22754 37214 22766 37266
rect 22818 37214 22830 37266
rect 24322 37214 24334 37266
rect 24386 37214 24398 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 27010 37214 27022 37266
rect 27074 37214 27086 37266
rect 31042 37214 31054 37266
rect 31106 37214 31118 37266
rect 19854 37202 19906 37214
rect 29262 37202 29314 37214
rect 31278 37202 31330 37214
rect 31502 37266 31554 37278
rect 31502 37202 31554 37214
rect 31614 37266 31666 37278
rect 31614 37202 31666 37214
rect 33742 37266 33794 37278
rect 33742 37202 33794 37214
rect 34190 37266 34242 37278
rect 34190 37202 34242 37214
rect 34414 37266 34466 37278
rect 34414 37202 34466 37214
rect 35198 37266 35250 37278
rect 39230 37266 39282 37278
rect 37986 37214 37998 37266
rect 38050 37214 38062 37266
rect 35198 37202 35250 37214
rect 39230 37202 39282 37214
rect 39566 37266 39618 37278
rect 43710 37266 43762 37278
rect 39778 37214 39790 37266
rect 39842 37214 39854 37266
rect 40898 37214 40910 37266
rect 40962 37214 40974 37266
rect 41794 37214 41806 37266
rect 41858 37214 41870 37266
rect 39566 37202 39618 37214
rect 43710 37202 43762 37214
rect 44382 37266 44434 37278
rect 44382 37202 44434 37214
rect 16830 37154 16882 37166
rect 28030 37154 28082 37166
rect 13682 37102 13694 37154
rect 13746 37102 13758 37154
rect 21522 37102 21534 37154
rect 21586 37102 21598 37154
rect 26338 37102 26350 37154
rect 26402 37102 26414 37154
rect 16830 37090 16882 37102
rect 28030 37090 28082 37102
rect 29822 37154 29874 37166
rect 29822 37090 29874 37102
rect 30270 37154 30322 37166
rect 30270 37090 30322 37102
rect 30718 37154 30770 37166
rect 30718 37090 30770 37102
rect 31390 37154 31442 37166
rect 31390 37090 31442 37102
rect 34750 37154 34802 37166
rect 40014 37154 40066 37166
rect 37762 37102 37774 37154
rect 37826 37102 37838 37154
rect 34750 37090 34802 37102
rect 40014 37090 40066 37102
rect 43822 37154 43874 37166
rect 43822 37090 43874 37102
rect 46958 37154 47010 37166
rect 46958 37090 47010 37102
rect 34974 37042 35026 37054
rect 12898 36990 12910 37042
rect 12962 36990 12974 37042
rect 14354 36990 14366 37042
rect 14418 36990 14430 37042
rect 34974 36978 35026 36990
rect 40126 37042 40178 37054
rect 40126 36978 40178 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 17614 36706 17666 36718
rect 44382 36706 44434 36718
rect 25106 36654 25118 36706
rect 25170 36654 25182 36706
rect 28466 36654 28478 36706
rect 28530 36654 28542 36706
rect 47394 36654 47406 36706
rect 47458 36654 47470 36706
rect 17614 36642 17666 36654
rect 44382 36642 44434 36654
rect 11230 36594 11282 36606
rect 18734 36594 18786 36606
rect 12450 36542 12462 36594
rect 12514 36542 12526 36594
rect 13794 36542 13806 36594
rect 13858 36542 13870 36594
rect 11230 36530 11282 36542
rect 18734 36530 18786 36542
rect 18958 36594 19010 36606
rect 34302 36594 34354 36606
rect 47070 36594 47122 36606
rect 20066 36542 20078 36594
rect 20130 36542 20142 36594
rect 26786 36542 26798 36594
rect 26850 36542 26862 36594
rect 29250 36542 29262 36594
rect 29314 36542 29326 36594
rect 30258 36542 30270 36594
rect 30322 36542 30334 36594
rect 39442 36542 39454 36594
rect 39506 36542 39518 36594
rect 45602 36542 45614 36594
rect 45666 36542 45678 36594
rect 18958 36530 19010 36542
rect 34302 36530 34354 36542
rect 47070 36530 47122 36542
rect 57934 36594 57986 36606
rect 57934 36530 57986 36542
rect 15822 36482 15874 36494
rect 18622 36482 18674 36494
rect 27918 36482 27970 36494
rect 10994 36430 11006 36482
rect 11058 36430 11070 36482
rect 14914 36430 14926 36482
rect 14978 36430 14990 36482
rect 16482 36430 16494 36482
rect 16546 36430 16558 36482
rect 16706 36430 16718 36482
rect 16770 36430 16782 36482
rect 17378 36430 17390 36482
rect 17442 36430 17454 36482
rect 19282 36430 19294 36482
rect 19346 36430 19358 36482
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 21522 36430 21534 36482
rect 21586 36430 21598 36482
rect 22754 36430 22766 36482
rect 22818 36430 22830 36482
rect 23538 36430 23550 36482
rect 23602 36430 23614 36482
rect 24546 36430 24558 36482
rect 24610 36430 24622 36482
rect 26002 36430 26014 36482
rect 26066 36430 26078 36482
rect 27122 36430 27134 36482
rect 27186 36430 27198 36482
rect 15822 36418 15874 36430
rect 18622 36418 18674 36430
rect 27918 36418 27970 36430
rect 28142 36482 28194 36494
rect 39118 36482 39170 36494
rect 42254 36482 42306 36494
rect 29138 36430 29150 36482
rect 29202 36430 29214 36482
rect 30594 36430 30606 36482
rect 30658 36430 30670 36482
rect 31042 36430 31054 36482
rect 31106 36430 31118 36482
rect 32386 36430 32398 36482
rect 32450 36430 32462 36482
rect 32722 36430 32734 36482
rect 32786 36430 32798 36482
rect 33058 36430 33070 36482
rect 33122 36430 33134 36482
rect 35634 36430 35646 36482
rect 35698 36430 35710 36482
rect 37874 36430 37886 36482
rect 37938 36430 37950 36482
rect 40898 36430 40910 36482
rect 40962 36430 40974 36482
rect 28142 36418 28194 36430
rect 39118 36418 39170 36430
rect 42254 36418 42306 36430
rect 42590 36482 42642 36494
rect 46846 36482 46898 36494
rect 42802 36430 42814 36482
rect 42866 36430 42878 36482
rect 44034 36430 44046 36482
rect 44098 36430 44110 36482
rect 45826 36430 45838 36482
rect 45890 36430 45902 36482
rect 55570 36430 55582 36482
rect 55634 36430 55646 36482
rect 42590 36418 42642 36430
rect 46846 36418 46898 36430
rect 9998 36370 10050 36382
rect 19518 36370 19570 36382
rect 41582 36370 41634 36382
rect 14018 36318 14030 36370
rect 14082 36318 14094 36370
rect 20738 36318 20750 36370
rect 20802 36318 20814 36370
rect 29250 36318 29262 36370
rect 29314 36318 29326 36370
rect 34514 36318 34526 36370
rect 34578 36318 34590 36370
rect 37986 36318 37998 36370
rect 38050 36318 38062 36370
rect 38770 36318 38782 36370
rect 38834 36318 38846 36370
rect 39890 36318 39902 36370
rect 39954 36318 39966 36370
rect 9998 36306 10050 36318
rect 19518 36306 19570 36318
rect 41582 36306 41634 36318
rect 41918 36370 41970 36382
rect 41918 36306 41970 36318
rect 42030 36370 42082 36382
rect 42030 36306 42082 36318
rect 43486 36370 43538 36382
rect 43486 36306 43538 36318
rect 43822 36370 43874 36382
rect 43822 36306 43874 36318
rect 46510 36370 46562 36382
rect 46510 36306 46562 36318
rect 9214 36258 9266 36270
rect 12910 36258 12962 36270
rect 11442 36206 11454 36258
rect 11506 36206 11518 36258
rect 9214 36194 9266 36206
rect 12910 36194 12962 36206
rect 44270 36258 44322 36270
rect 44270 36194 44322 36206
rect 44830 36258 44882 36270
rect 45154 36206 45166 36258
rect 45218 36206 45230 36258
rect 44830 36194 44882 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 24222 35922 24274 35934
rect 13234 35870 13246 35922
rect 13298 35870 13310 35922
rect 14578 35870 14590 35922
rect 14642 35870 14654 35922
rect 23538 35870 23550 35922
rect 23602 35870 23614 35922
rect 24222 35858 24274 35870
rect 24446 35922 24498 35934
rect 30606 35922 30658 35934
rect 29026 35870 29038 35922
rect 29090 35870 29102 35922
rect 24446 35858 24498 35870
rect 30606 35858 30658 35870
rect 32174 35922 32226 35934
rect 34862 35922 34914 35934
rect 34178 35870 34190 35922
rect 34242 35870 34254 35922
rect 32174 35858 32226 35870
rect 34862 35858 34914 35870
rect 35534 35922 35586 35934
rect 35534 35858 35586 35870
rect 35646 35922 35698 35934
rect 35646 35858 35698 35870
rect 36878 35922 36930 35934
rect 40014 35922 40066 35934
rect 39666 35870 39678 35922
rect 39730 35870 39742 35922
rect 36878 35858 36930 35870
rect 40014 35858 40066 35870
rect 42702 35922 42754 35934
rect 43026 35870 43038 35922
rect 43090 35870 43102 35922
rect 42702 35858 42754 35870
rect 9550 35810 9602 35822
rect 7858 35758 7870 35810
rect 7922 35758 7934 35810
rect 9550 35746 9602 35758
rect 11342 35810 11394 35822
rect 15710 35810 15762 35822
rect 31726 35810 31778 35822
rect 11666 35758 11678 35810
rect 11730 35758 11742 35810
rect 14130 35758 14142 35810
rect 14194 35758 14206 35810
rect 27570 35758 27582 35810
rect 27634 35758 27646 35810
rect 30146 35758 30158 35810
rect 30210 35758 30222 35810
rect 11342 35746 11394 35758
rect 15710 35746 15762 35758
rect 31726 35746 31778 35758
rect 34526 35810 34578 35822
rect 34526 35746 34578 35758
rect 34638 35810 34690 35822
rect 34638 35746 34690 35758
rect 44494 35810 44546 35822
rect 46722 35758 46734 35810
rect 46786 35758 46798 35810
rect 44494 35746 44546 35758
rect 10782 35698 10834 35710
rect 16046 35698 16098 35710
rect 8754 35646 8766 35698
rect 8818 35646 8830 35698
rect 9986 35646 9998 35698
rect 10050 35646 10062 35698
rect 11890 35646 11902 35698
rect 11954 35646 11966 35698
rect 13682 35646 13694 35698
rect 13746 35646 13758 35698
rect 14578 35646 14590 35698
rect 14642 35646 14654 35698
rect 15250 35646 15262 35698
rect 15314 35646 15326 35698
rect 10782 35634 10834 35646
rect 16046 35634 16098 35646
rect 17726 35698 17778 35710
rect 23214 35698 23266 35710
rect 18498 35646 18510 35698
rect 18562 35646 18574 35698
rect 19394 35646 19406 35698
rect 19458 35646 19470 35698
rect 20962 35646 20974 35698
rect 21026 35646 21038 35698
rect 21410 35646 21422 35698
rect 21474 35646 21486 35698
rect 17726 35634 17778 35646
rect 23214 35634 23266 35646
rect 24670 35698 24722 35710
rect 30942 35698 30994 35710
rect 25330 35646 25342 35698
rect 25394 35646 25406 35698
rect 25554 35646 25566 35698
rect 25618 35646 25630 35698
rect 26674 35646 26686 35698
rect 26738 35646 26750 35698
rect 27458 35646 27470 35698
rect 27522 35646 27534 35698
rect 28914 35646 28926 35698
rect 28978 35646 28990 35698
rect 24670 35634 24722 35646
rect 30942 35634 30994 35646
rect 33854 35698 33906 35710
rect 33854 35634 33906 35646
rect 34974 35698 35026 35710
rect 34974 35634 35026 35646
rect 35422 35698 35474 35710
rect 35422 35634 35474 35646
rect 36206 35698 36258 35710
rect 36206 35634 36258 35646
rect 36430 35698 36482 35710
rect 36430 35634 36482 35646
rect 43598 35698 43650 35710
rect 43922 35646 43934 35698
rect 43986 35646 43998 35698
rect 46498 35646 46510 35698
rect 46562 35646 46574 35698
rect 43598 35634 43650 35646
rect 16606 35586 16658 35598
rect 16606 35522 16658 35534
rect 17502 35586 17554 35598
rect 24558 35586 24610 35598
rect 33630 35586 33682 35598
rect 18050 35534 18062 35586
rect 18114 35534 18126 35586
rect 21858 35534 21870 35586
rect 21922 35534 21934 35586
rect 26226 35534 26238 35586
rect 26290 35534 26302 35586
rect 30594 35534 30606 35586
rect 30658 35534 30670 35586
rect 17502 35522 17554 35534
rect 24558 35522 24610 35534
rect 33630 35522 33682 35534
rect 35982 35586 36034 35598
rect 35982 35522 36034 35534
rect 21746 35422 21758 35474
rect 21810 35422 21822 35474
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 19406 35138 19458 35150
rect 9314 35086 9326 35138
rect 9378 35086 9390 35138
rect 17378 35086 17390 35138
rect 17442 35086 17454 35138
rect 19406 35074 19458 35086
rect 25006 35138 25058 35150
rect 25006 35074 25058 35086
rect 28590 35138 28642 35150
rect 28590 35074 28642 35086
rect 29822 35138 29874 35150
rect 29822 35074 29874 35086
rect 31166 35138 31218 35150
rect 31166 35074 31218 35086
rect 15374 35026 15426 35038
rect 19966 35026 20018 35038
rect 24894 35026 24946 35038
rect 28142 35026 28194 35038
rect 32398 35026 32450 35038
rect 10770 34974 10782 35026
rect 10834 34974 10846 35026
rect 14018 34974 14030 35026
rect 14082 34974 14094 35026
rect 18386 34974 18398 35026
rect 18450 34974 18462 35026
rect 21746 34974 21758 35026
rect 21810 34974 21822 35026
rect 24210 34974 24222 35026
rect 24274 34974 24286 35026
rect 27346 34974 27358 35026
rect 27410 34974 27422 35026
rect 30258 34974 30270 35026
rect 30322 34974 30334 35026
rect 15374 34962 15426 34974
rect 19966 34962 20018 34974
rect 24894 34962 24946 34974
rect 28142 34962 28194 34974
rect 32398 34962 32450 34974
rect 34638 35026 34690 35038
rect 34638 34962 34690 34974
rect 36318 35026 36370 35038
rect 40674 34974 40686 35026
rect 40738 34974 40750 35026
rect 57810 34974 57822 35026
rect 57874 34974 57886 35026
rect 36318 34962 36370 34974
rect 8766 34914 8818 34926
rect 8766 34850 8818 34862
rect 8990 34914 9042 34926
rect 14814 34914 14866 34926
rect 25790 34914 25842 34926
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 11778 34862 11790 34914
rect 11842 34862 11854 34914
rect 12898 34862 12910 34914
rect 12962 34862 12974 34914
rect 16034 34862 16046 34914
rect 16098 34862 16110 34914
rect 19282 34862 19294 34914
rect 19346 34862 19358 34914
rect 23538 34862 23550 34914
rect 23602 34862 23614 34914
rect 8990 34850 9042 34862
rect 14814 34850 14866 34862
rect 25790 34850 25842 34862
rect 26014 34914 26066 34926
rect 29486 34914 29538 34926
rect 26674 34862 26686 34914
rect 26738 34862 26750 34914
rect 29250 34862 29262 34914
rect 29314 34862 29326 34914
rect 26014 34850 26066 34862
rect 29486 34850 29538 34862
rect 29710 34914 29762 34926
rect 35870 34914 35922 34926
rect 30594 34862 30606 34914
rect 30658 34862 30670 34914
rect 35074 34862 35086 34914
rect 35138 34862 35150 34914
rect 40338 34862 40350 34914
rect 40402 34862 40414 34914
rect 55570 34862 55582 34914
rect 55634 34862 55646 34914
rect 29710 34850 29762 34862
rect 35870 34850 35922 34862
rect 28478 34802 28530 34814
rect 16482 34750 16494 34802
rect 16546 34750 16558 34802
rect 19170 34750 19182 34802
rect 19234 34750 19246 34802
rect 20402 34750 20414 34802
rect 20466 34750 20478 34802
rect 22754 34750 22766 34802
rect 22818 34750 22830 34802
rect 27010 34750 27022 34802
rect 27074 34750 27086 34802
rect 28478 34738 28530 34750
rect 31054 34802 31106 34814
rect 31054 34738 31106 34750
rect 31166 34802 31218 34814
rect 31166 34738 31218 34750
rect 32510 34802 32562 34814
rect 32510 34738 32562 34750
rect 35534 34802 35586 34814
rect 41358 34802 41410 34814
rect 40002 34750 40014 34802
rect 40066 34750 40078 34802
rect 35534 34738 35586 34750
rect 41358 34738 41410 34750
rect 13582 34690 13634 34702
rect 13582 34626 13634 34638
rect 14478 34690 14530 34702
rect 14478 34626 14530 34638
rect 17950 34690 18002 34702
rect 17950 34626 18002 34638
rect 20750 34690 20802 34702
rect 20750 34626 20802 34638
rect 21310 34690 21362 34702
rect 21310 34626 21362 34638
rect 22318 34690 22370 34702
rect 22318 34626 22370 34638
rect 25454 34690 25506 34702
rect 41022 34690 41074 34702
rect 26338 34638 26350 34690
rect 26402 34638 26414 34690
rect 34850 34638 34862 34690
rect 34914 34638 34926 34690
rect 25454 34626 25506 34638
rect 41022 34626 41074 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 14926 34354 14978 34366
rect 16830 34354 16882 34366
rect 15698 34302 15710 34354
rect 15762 34302 15774 34354
rect 14926 34290 14978 34302
rect 16830 34290 16882 34302
rect 17726 34354 17778 34366
rect 33406 34354 33458 34366
rect 19170 34302 19182 34354
rect 19234 34302 19246 34354
rect 17726 34290 17778 34302
rect 33406 34290 33458 34302
rect 33854 34354 33906 34366
rect 33854 34290 33906 34302
rect 38110 34354 38162 34366
rect 43374 34354 43426 34366
rect 41458 34302 41470 34354
rect 41522 34302 41534 34354
rect 38110 34290 38162 34302
rect 43374 34290 43426 34302
rect 44494 34354 44546 34366
rect 44494 34290 44546 34302
rect 14702 34242 14754 34254
rect 24334 34242 24386 34254
rect 10658 34190 10670 34242
rect 10722 34190 10734 34242
rect 19842 34190 19854 34242
rect 19906 34190 19918 34242
rect 14702 34178 14754 34190
rect 24334 34178 24386 34190
rect 24446 34242 24498 34254
rect 24446 34178 24498 34190
rect 24670 34242 24722 34254
rect 37326 34242 37378 34254
rect 31826 34190 31838 34242
rect 31890 34190 31902 34242
rect 33058 34190 33070 34242
rect 33122 34190 33134 34242
rect 24670 34178 24722 34190
rect 37326 34178 37378 34190
rect 58158 34242 58210 34254
rect 58158 34178 58210 34190
rect 8990 34130 9042 34142
rect 10110 34130 10162 34142
rect 14590 34130 14642 34142
rect 4162 34078 4174 34130
rect 4226 34078 4238 34130
rect 9650 34078 9662 34130
rect 9714 34078 9726 34130
rect 11106 34078 11118 34130
rect 11170 34078 11182 34130
rect 12338 34078 12350 34130
rect 12402 34078 12414 34130
rect 13570 34078 13582 34130
rect 13634 34078 13646 34130
rect 8990 34066 9042 34078
rect 10110 34066 10162 34078
rect 14590 34066 14642 34078
rect 16270 34130 16322 34142
rect 16270 34066 16322 34078
rect 18286 34130 18338 34142
rect 18286 34066 18338 34078
rect 18622 34130 18674 34142
rect 18622 34066 18674 34078
rect 18846 34130 18898 34142
rect 30718 34130 30770 34142
rect 20178 34078 20190 34130
rect 20242 34078 20254 34130
rect 22642 34078 22654 34130
rect 22706 34078 22718 34130
rect 23202 34078 23214 34130
rect 23266 34078 23278 34130
rect 26114 34078 26126 34130
rect 26178 34078 26190 34130
rect 28354 34078 28366 34130
rect 28418 34078 28430 34130
rect 28690 34078 28702 34130
rect 28754 34078 28766 34130
rect 29026 34078 29038 34130
rect 29090 34078 29102 34130
rect 18846 34066 18898 34078
rect 30718 34066 30770 34078
rect 32174 34130 32226 34142
rect 32174 34066 32226 34078
rect 34414 34130 34466 34142
rect 39790 34130 39842 34142
rect 34962 34078 34974 34130
rect 35026 34078 35038 34130
rect 39106 34078 39118 34130
rect 39170 34078 39182 34130
rect 34414 34066 34466 34078
rect 39790 34066 39842 34078
rect 40910 34130 40962 34142
rect 40910 34066 40962 34078
rect 41134 34130 41186 34142
rect 41134 34066 41186 34078
rect 43150 34130 43202 34142
rect 43150 34066 43202 34078
rect 43486 34130 43538 34142
rect 43486 34066 43538 34078
rect 44158 34130 44210 34142
rect 44158 34066 44210 34078
rect 44606 34130 44658 34142
rect 44606 34066 44658 34078
rect 4846 34018 4898 34030
rect 15150 34018 15202 34030
rect 25566 34018 25618 34030
rect 8530 33966 8542 34018
rect 8594 33966 8606 34018
rect 11666 33966 11678 34018
rect 11730 33966 11742 34018
rect 20962 33966 20974 34018
rect 21026 33966 21038 34018
rect 26562 33966 26574 34018
rect 26626 33966 26638 34018
rect 31154 33966 31166 34018
rect 31218 33966 31230 34018
rect 39442 33966 39454 34018
rect 39506 33966 39518 34018
rect 4846 33954 4898 33966
rect 15150 33954 15202 33966
rect 25566 33954 25618 33966
rect 1934 33906 1986 33918
rect 1934 33842 1986 33854
rect 15374 33906 15426 33918
rect 15374 33842 15426 33854
rect 23886 33906 23938 33918
rect 23886 33842 23938 33854
rect 24110 33906 24162 33918
rect 30034 33854 30046 33906
rect 30098 33854 30110 33906
rect 24110 33842 24162 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 10446 33570 10498 33582
rect 10446 33506 10498 33518
rect 19518 33570 19570 33582
rect 19518 33506 19570 33518
rect 25678 33570 25730 33582
rect 25678 33506 25730 33518
rect 35198 33570 35250 33582
rect 38098 33567 38110 33570
rect 35198 33506 35250 33518
rect 37777 33521 38110 33567
rect 1934 33458 1986 33470
rect 14814 33458 14866 33470
rect 12226 33406 12238 33458
rect 12290 33406 12302 33458
rect 1934 33394 1986 33406
rect 14814 33394 14866 33406
rect 17838 33458 17890 33470
rect 17838 33394 17890 33406
rect 18062 33458 18114 33470
rect 24670 33458 24722 33470
rect 18610 33406 18622 33458
rect 18674 33406 18686 33458
rect 19282 33406 19294 33458
rect 19346 33406 19358 33458
rect 20290 33406 20302 33458
rect 20354 33406 20366 33458
rect 23202 33406 23214 33458
rect 23266 33406 23278 33458
rect 18062 33394 18114 33406
rect 24670 33394 24722 33406
rect 25342 33458 25394 33470
rect 26798 33458 26850 33470
rect 26226 33406 26238 33458
rect 26290 33406 26302 33458
rect 25342 33394 25394 33406
rect 26798 33394 26850 33406
rect 27134 33458 27186 33470
rect 29822 33458 29874 33470
rect 37777 33458 37823 33521
rect 38098 33518 38110 33521
rect 38162 33518 38174 33570
rect 28130 33406 28142 33458
rect 28194 33406 28206 33458
rect 37426 33406 37438 33458
rect 37490 33406 37502 33458
rect 37762 33406 37774 33458
rect 37826 33406 37838 33458
rect 27134 33394 27186 33406
rect 29822 33394 29874 33406
rect 9998 33346 10050 33358
rect 4274 33294 4286 33346
rect 4338 33294 4350 33346
rect 9998 33282 10050 33294
rect 10558 33346 10610 33358
rect 10558 33282 10610 33294
rect 10782 33346 10834 33358
rect 24222 33346 24274 33358
rect 12674 33294 12686 33346
rect 12738 33294 12750 33346
rect 16594 33294 16606 33346
rect 16658 33294 16670 33346
rect 17042 33294 17054 33346
rect 17106 33294 17118 33346
rect 18498 33294 18510 33346
rect 18562 33294 18574 33346
rect 22082 33294 22094 33346
rect 22146 33294 22158 33346
rect 22642 33294 22654 33346
rect 22706 33294 22718 33346
rect 23426 33294 23438 33346
rect 23490 33294 23502 33346
rect 10782 33282 10834 33294
rect 24222 33282 24274 33294
rect 25454 33346 25506 33358
rect 30382 33346 30434 33358
rect 31502 33346 31554 33358
rect 35646 33346 35698 33358
rect 27570 33294 27582 33346
rect 27634 33294 27646 33346
rect 28466 33294 28478 33346
rect 28530 33294 28542 33346
rect 29362 33294 29374 33346
rect 29426 33294 29438 33346
rect 30930 33294 30942 33346
rect 30994 33294 31006 33346
rect 32162 33294 32174 33346
rect 32226 33294 32238 33346
rect 25454 33282 25506 33294
rect 30382 33282 30434 33294
rect 31502 33282 31554 33294
rect 35646 33282 35698 33294
rect 36990 33346 37042 33358
rect 36990 33282 37042 33294
rect 40014 33346 40066 33358
rect 43038 33346 43090 33358
rect 42130 33294 42142 33346
rect 42194 33294 42206 33346
rect 45042 33294 45054 33346
rect 45106 33294 45118 33346
rect 40014 33282 40066 33294
rect 43038 33282 43090 33294
rect 15598 33234 15650 33246
rect 24558 33234 24610 33246
rect 30718 33234 30770 33246
rect 17266 33182 17278 33234
rect 17330 33182 17342 33234
rect 29138 33182 29150 33234
rect 29202 33182 29214 33234
rect 15598 33170 15650 33182
rect 24558 33170 24610 33182
rect 30718 33170 30770 33182
rect 40350 33234 40402 33246
rect 40350 33170 40402 33182
rect 42926 33234 42978 33246
rect 42926 33170 42978 33182
rect 9438 33122 9490 33134
rect 9438 33058 9490 33070
rect 11230 33122 11282 33134
rect 11230 33058 11282 33070
rect 16494 33122 16546 33134
rect 16494 33058 16546 33070
rect 19294 33122 19346 33134
rect 19294 33058 19346 33070
rect 20750 33122 20802 33134
rect 20750 33058 20802 33070
rect 21758 33122 21810 33134
rect 21758 33058 21810 33070
rect 23662 33122 23714 33134
rect 23662 33058 23714 33070
rect 24782 33122 24834 33134
rect 37998 33122 38050 33134
rect 34402 33070 34414 33122
rect 34466 33070 34478 33122
rect 24782 33058 24834 33070
rect 37998 33058 38050 33070
rect 38782 33122 38834 33134
rect 38782 33058 38834 33070
rect 41918 33122 41970 33134
rect 41918 33058 41970 33070
rect 42702 33122 42754 33134
rect 42702 33058 42754 33070
rect 44830 33122 44882 33134
rect 44830 33058 44882 33070
rect 58158 33122 58210 33134
rect 58158 33058 58210 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 13470 32786 13522 32798
rect 13470 32722 13522 32734
rect 15934 32786 15986 32798
rect 15934 32722 15986 32734
rect 20750 32786 20802 32798
rect 20750 32722 20802 32734
rect 22430 32786 22482 32798
rect 25902 32786 25954 32798
rect 23874 32734 23886 32786
rect 23938 32734 23950 32786
rect 22430 32722 22482 32734
rect 25902 32722 25954 32734
rect 27918 32786 27970 32798
rect 27918 32722 27970 32734
rect 28702 32786 28754 32798
rect 29374 32786 29426 32798
rect 29026 32734 29038 32786
rect 29090 32734 29102 32786
rect 28702 32722 28754 32734
rect 29374 32722 29426 32734
rect 29710 32786 29762 32798
rect 29710 32722 29762 32734
rect 30382 32786 30434 32798
rect 30382 32722 30434 32734
rect 37438 32786 37490 32798
rect 37438 32722 37490 32734
rect 38110 32786 38162 32798
rect 38110 32722 38162 32734
rect 39454 32786 39506 32798
rect 39454 32722 39506 32734
rect 39678 32786 39730 32798
rect 39678 32722 39730 32734
rect 45390 32786 45442 32798
rect 45390 32722 45442 32734
rect 1710 32674 1762 32686
rect 1710 32610 1762 32622
rect 8878 32674 8930 32686
rect 8878 32610 8930 32622
rect 13582 32674 13634 32686
rect 15710 32674 15762 32686
rect 22878 32674 22930 32686
rect 14242 32622 14254 32674
rect 14306 32622 14318 32674
rect 19058 32622 19070 32674
rect 19122 32622 19134 32674
rect 13582 32610 13634 32622
rect 15710 32610 15762 32622
rect 22878 32610 22930 32622
rect 24670 32674 24722 32686
rect 36878 32674 36930 32686
rect 31602 32622 31614 32674
rect 31666 32622 31678 32674
rect 24670 32610 24722 32622
rect 36878 32610 36930 32622
rect 37214 32674 37266 32686
rect 37214 32610 37266 32622
rect 38334 32674 38386 32686
rect 38334 32610 38386 32622
rect 39118 32674 39170 32686
rect 39118 32610 39170 32622
rect 44606 32674 44658 32686
rect 44606 32610 44658 32622
rect 9774 32562 9826 32574
rect 9774 32498 9826 32510
rect 10670 32562 10722 32574
rect 10670 32498 10722 32510
rect 11230 32562 11282 32574
rect 14814 32562 14866 32574
rect 12450 32510 12462 32562
rect 12514 32510 12526 32562
rect 14018 32510 14030 32562
rect 14082 32510 14094 32562
rect 11230 32498 11282 32510
rect 14814 32498 14866 32510
rect 15598 32562 15650 32574
rect 19406 32562 19458 32574
rect 17826 32510 17838 32562
rect 17890 32510 17902 32562
rect 15598 32498 15650 32510
rect 19406 32498 19458 32510
rect 19966 32562 20018 32574
rect 25454 32562 25506 32574
rect 37886 32562 37938 32574
rect 21410 32510 21422 32562
rect 21474 32510 21486 32562
rect 21634 32510 21646 32562
rect 21698 32510 21710 32562
rect 23314 32510 23326 32562
rect 23378 32510 23390 32562
rect 24098 32510 24110 32562
rect 24162 32510 24174 32562
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 19966 32498 20018 32510
rect 25454 32498 25506 32510
rect 37886 32498 37938 32510
rect 38222 32562 38274 32574
rect 38222 32498 38274 32510
rect 38782 32562 38834 32574
rect 38782 32498 38834 32510
rect 38894 32562 38946 32574
rect 38894 32498 38946 32510
rect 39230 32562 39282 32574
rect 39230 32498 39282 32510
rect 39790 32562 39842 32574
rect 39790 32498 39842 32510
rect 41694 32562 41746 32574
rect 42242 32510 42254 32562
rect 42306 32510 42318 32562
rect 41694 32498 41746 32510
rect 15150 32450 15202 32462
rect 29822 32450 29874 32462
rect 10210 32398 10222 32450
rect 10274 32398 10286 32450
rect 12114 32398 12126 32450
rect 12178 32398 12190 32450
rect 17938 32398 17950 32450
rect 18002 32398 18014 32450
rect 21522 32398 21534 32450
rect 21586 32398 21598 32450
rect 15150 32386 15202 32398
rect 29822 32386 29874 32398
rect 37326 32450 37378 32462
rect 37326 32386 37378 32398
rect 8990 32338 9042 32350
rect 8990 32274 9042 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 24446 32002 24498 32014
rect 24446 31938 24498 31950
rect 40126 32002 40178 32014
rect 40126 31938 40178 31950
rect 1934 31890 1986 31902
rect 1934 31826 1986 31838
rect 10558 31890 10610 31902
rect 10558 31826 10610 31838
rect 11454 31890 11506 31902
rect 11454 31826 11506 31838
rect 14702 31890 14754 31902
rect 14702 31826 14754 31838
rect 18846 31890 18898 31902
rect 18846 31826 18898 31838
rect 21758 31890 21810 31902
rect 21758 31826 21810 31838
rect 22542 31890 22594 31902
rect 22542 31826 22594 31838
rect 23998 31890 24050 31902
rect 23998 31826 24050 31838
rect 29374 31890 29426 31902
rect 29374 31826 29426 31838
rect 9998 31778 10050 31790
rect 4274 31726 4286 31778
rect 4338 31726 4350 31778
rect 9998 31714 10050 31726
rect 10894 31778 10946 31790
rect 10894 31714 10946 31726
rect 11790 31778 11842 31790
rect 11790 31714 11842 31726
rect 14142 31778 14194 31790
rect 14142 31714 14194 31726
rect 21982 31666 22034 31678
rect 24334 31666 24386 31678
rect 12114 31614 12126 31666
rect 12178 31614 12190 31666
rect 23202 31614 23214 31666
rect 23266 31614 23278 31666
rect 21982 31602 22034 31614
rect 24334 31602 24386 31614
rect 25454 31666 25506 31678
rect 38210 31614 38222 31666
rect 38274 31614 38286 31666
rect 25454 31602 25506 31614
rect 4734 31554 4786 31566
rect 4734 31490 4786 31502
rect 22878 31554 22930 31566
rect 22878 31490 22930 31502
rect 24446 31554 24498 31566
rect 24446 31490 24498 31502
rect 25006 31554 25058 31566
rect 25006 31490 25058 31502
rect 25566 31554 25618 31566
rect 25566 31490 25618 31502
rect 25790 31554 25842 31566
rect 25790 31490 25842 31502
rect 26462 31554 26514 31566
rect 26462 31490 26514 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 9102 31218 9154 31230
rect 18286 31218 18338 31230
rect 19742 31218 19794 31230
rect 8530 31166 8542 31218
rect 8594 31166 8606 31218
rect 12338 31166 12350 31218
rect 12402 31166 12414 31218
rect 13346 31166 13358 31218
rect 13410 31166 13422 31218
rect 14466 31166 14478 31218
rect 14530 31166 14542 31218
rect 18946 31166 18958 31218
rect 19010 31166 19022 31218
rect 9102 31154 9154 31166
rect 18286 31154 18338 31166
rect 19742 31154 19794 31166
rect 20302 31218 20354 31230
rect 20302 31154 20354 31166
rect 22206 31218 22258 31230
rect 22206 31154 22258 31166
rect 23438 31218 23490 31230
rect 23438 31154 23490 31166
rect 23550 31218 23602 31230
rect 23550 31154 23602 31166
rect 23774 31218 23826 31230
rect 23774 31154 23826 31166
rect 24446 31218 24498 31230
rect 24446 31154 24498 31166
rect 24670 31218 24722 31230
rect 24670 31154 24722 31166
rect 30158 31218 30210 31230
rect 45278 31218 45330 31230
rect 44594 31166 44606 31218
rect 44658 31166 44670 31218
rect 30158 31154 30210 31166
rect 45278 31154 45330 31166
rect 9550 31106 9602 31118
rect 19630 31106 19682 31118
rect 16706 31054 16718 31106
rect 16770 31054 16782 31106
rect 9550 31042 9602 31054
rect 19630 31042 19682 31054
rect 23886 31106 23938 31118
rect 23886 31042 23938 31054
rect 29374 31106 29426 31118
rect 29374 31042 29426 31054
rect 35870 31106 35922 31118
rect 57822 31106 57874 31118
rect 38882 31054 38894 31106
rect 38946 31054 38958 31106
rect 35870 31042 35922 31054
rect 57822 31042 57874 31054
rect 5630 30994 5682 31006
rect 13022 30994 13074 31006
rect 4274 30942 4286 30994
rect 4338 30942 4350 30994
rect 6066 30942 6078 30994
rect 6130 30942 6142 30994
rect 9762 30942 9774 30994
rect 9826 30942 9838 30994
rect 12562 30942 12574 30994
rect 12626 30942 12638 30994
rect 5630 30930 5682 30942
rect 13022 30930 13074 30942
rect 14814 30994 14866 31006
rect 18062 30994 18114 31006
rect 15810 30942 15822 30994
rect 15874 30942 15886 30994
rect 14814 30930 14866 30942
rect 18062 30930 18114 30942
rect 18174 30994 18226 31006
rect 18174 30930 18226 30942
rect 18734 30994 18786 31006
rect 21310 30994 21362 31006
rect 32958 30994 33010 31006
rect 58158 30994 58210 31006
rect 19170 30942 19182 30994
rect 19234 30942 19246 30994
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 24210 30942 24222 30994
rect 24274 30942 24286 30994
rect 25778 30942 25790 30994
rect 25842 30942 25854 30994
rect 26562 30942 26574 30994
rect 26626 30942 26638 30994
rect 27010 30942 27022 30994
rect 27074 30942 27086 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 38658 30942 38670 30994
rect 38722 30942 38734 30994
rect 41682 30942 41694 30994
rect 41746 30942 41758 30994
rect 42242 30942 42254 30994
rect 42306 30942 42318 30994
rect 18734 30930 18786 30942
rect 21310 30930 21362 30942
rect 32958 30930 33010 30942
rect 58158 30930 58210 30942
rect 1934 30882 1986 30894
rect 20974 30882 21026 30894
rect 15698 30830 15710 30882
rect 15762 30830 15774 30882
rect 1934 30818 1986 30830
rect 20974 30818 21026 30830
rect 22318 30882 22370 30894
rect 22318 30818 22370 30830
rect 22766 30882 22818 30894
rect 26238 30882 26290 30894
rect 24658 30830 24670 30882
rect 24722 30830 24734 30882
rect 25330 30830 25342 30882
rect 25394 30830 25406 30882
rect 22766 30818 22818 30830
rect 26238 30818 26290 30830
rect 57598 30882 57650 30894
rect 57598 30818 57650 30830
rect 19742 30770 19794 30782
rect 19742 30706 19794 30718
rect 36654 30770 36706 30782
rect 36654 30706 36706 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 25342 30434 25394 30446
rect 16594 30382 16606 30434
rect 16658 30382 16670 30434
rect 25342 30370 25394 30382
rect 26462 30434 26514 30446
rect 26462 30370 26514 30382
rect 26798 30434 26850 30446
rect 26798 30370 26850 30382
rect 38894 30434 38946 30446
rect 38894 30370 38946 30382
rect 1710 30322 1762 30334
rect 1710 30258 1762 30270
rect 21870 30322 21922 30334
rect 23874 30270 23886 30322
rect 23938 30270 23950 30322
rect 36194 30270 36206 30322
rect 36258 30270 36270 30322
rect 21870 30258 21922 30270
rect 9102 30210 9154 30222
rect 12574 30210 12626 30222
rect 16494 30210 16546 30222
rect 12226 30158 12238 30210
rect 12290 30158 12302 30210
rect 15810 30158 15822 30210
rect 15874 30158 15886 30210
rect 9102 30146 9154 30158
rect 12574 30146 12626 30158
rect 16494 30146 16546 30158
rect 17390 30210 17442 30222
rect 17390 30146 17442 30158
rect 17838 30210 17890 30222
rect 17838 30146 17890 30158
rect 17950 30210 18002 30222
rect 17950 30146 18002 30158
rect 18622 30210 18674 30222
rect 29822 30210 29874 30222
rect 33294 30210 33346 30222
rect 23650 30158 23662 30210
rect 23714 30158 23726 30210
rect 30258 30158 30270 30210
rect 30322 30158 30334 30210
rect 18622 30146 18674 30158
rect 29822 30146 29874 30158
rect 33294 30146 33346 30158
rect 34750 30210 34802 30222
rect 35522 30158 35534 30210
rect 35586 30158 35598 30210
rect 34750 30146 34802 30158
rect 17726 30098 17778 30110
rect 17726 30034 17778 30046
rect 18286 30098 18338 30110
rect 18286 30034 18338 30046
rect 18734 30098 18786 30110
rect 18734 30034 18786 30046
rect 18958 30098 19010 30110
rect 18958 30034 19010 30046
rect 19182 30098 19234 30110
rect 19182 30034 19234 30046
rect 19630 30098 19682 30110
rect 19630 30034 19682 30046
rect 22990 30098 23042 30110
rect 22990 30034 23042 30046
rect 24334 30098 24386 30110
rect 24334 30034 24386 30046
rect 24558 30098 24610 30110
rect 24558 30034 24610 30046
rect 25790 30098 25842 30110
rect 25790 30034 25842 30046
rect 34862 30098 34914 30110
rect 35858 30046 35870 30098
rect 35922 30046 35934 30098
rect 34862 30034 34914 30046
rect 2158 29986 2210 29998
rect 15262 29986 15314 29998
rect 9650 29934 9662 29986
rect 9714 29934 9726 29986
rect 14914 29934 14926 29986
rect 14978 29934 14990 29986
rect 2158 29922 2210 29934
rect 15262 29922 15314 29934
rect 24446 29986 24498 29998
rect 24446 29922 24498 29934
rect 25118 29986 25170 29998
rect 25118 29922 25170 29934
rect 25230 29986 25282 29998
rect 25230 29922 25282 29934
rect 26686 29986 26738 29998
rect 34526 29986 34578 29998
rect 32722 29934 32734 29986
rect 32786 29934 32798 29986
rect 26686 29922 26738 29934
rect 34526 29922 34578 29934
rect 39118 29986 39170 29998
rect 39118 29922 39170 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 11790 29650 11842 29662
rect 23886 29650 23938 29662
rect 19618 29598 19630 29650
rect 19682 29598 19694 29650
rect 11790 29586 11842 29598
rect 23886 29586 23938 29598
rect 24670 29650 24722 29662
rect 24670 29586 24722 29598
rect 25454 29650 25506 29662
rect 25454 29586 25506 29598
rect 28590 29650 28642 29662
rect 28590 29586 28642 29598
rect 29822 29650 29874 29662
rect 39118 29650 39170 29662
rect 38098 29598 38110 29650
rect 38162 29598 38174 29650
rect 29822 29586 29874 29598
rect 39118 29586 39170 29598
rect 39566 29650 39618 29662
rect 39566 29586 39618 29598
rect 33406 29538 33458 29550
rect 33406 29474 33458 29486
rect 44494 29538 44546 29550
rect 44494 29474 44546 29486
rect 22542 29426 22594 29438
rect 34974 29426 35026 29438
rect 38894 29426 38946 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 12338 29374 12350 29426
rect 12402 29374 12414 29426
rect 22082 29374 22094 29426
rect 22146 29374 22158 29426
rect 24098 29374 24110 29426
rect 24162 29374 24174 29426
rect 28354 29374 28366 29426
rect 28418 29374 28430 29426
rect 30034 29374 30046 29426
rect 30098 29374 30110 29426
rect 33618 29374 33630 29426
rect 33682 29374 33694 29426
rect 35634 29374 35646 29426
rect 35698 29374 35710 29426
rect 22542 29362 22594 29374
rect 34974 29362 35026 29374
rect 38894 29362 38946 29374
rect 41582 29426 41634 29438
rect 42242 29374 42254 29426
rect 42306 29374 42318 29426
rect 41582 29362 41634 29374
rect 13022 29314 13074 29326
rect 12562 29262 12574 29314
rect 12626 29262 12638 29314
rect 13022 29250 13074 29262
rect 18958 29314 19010 29326
rect 18958 29250 19010 29262
rect 27918 29314 27970 29326
rect 27918 29250 27970 29262
rect 39678 29314 39730 29326
rect 39678 29250 39730 29262
rect 1934 29202 1986 29214
rect 1934 29138 1986 29150
rect 19070 29202 19122 29214
rect 19070 29138 19122 29150
rect 23774 29202 23826 29214
rect 23774 29138 23826 29150
rect 38670 29202 38722 29214
rect 38670 29138 38722 29150
rect 45278 29202 45330 29214
rect 45278 29138 45330 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 17054 28866 17106 28878
rect 17054 28802 17106 28814
rect 28478 28866 28530 28878
rect 28478 28802 28530 28814
rect 24446 28754 24498 28766
rect 24446 28690 24498 28702
rect 34302 28754 34354 28766
rect 34302 28690 34354 28702
rect 6302 28642 6354 28654
rect 25006 28642 25058 28654
rect 29150 28642 29202 28654
rect 12674 28590 12686 28642
rect 12738 28590 12750 28642
rect 13458 28590 13470 28642
rect 13522 28590 13534 28642
rect 13906 28590 13918 28642
rect 13970 28590 13982 28642
rect 20402 28590 20414 28642
rect 20466 28590 20478 28642
rect 25330 28590 25342 28642
rect 25394 28590 25406 28642
rect 6302 28578 6354 28590
rect 25006 28578 25058 28590
rect 29150 28578 29202 28590
rect 30046 28642 30098 28654
rect 33518 28642 33570 28654
rect 30370 28590 30382 28642
rect 30434 28590 30446 28642
rect 30046 28578 30098 28590
rect 33518 28578 33570 28590
rect 34078 28642 34130 28654
rect 34078 28578 34130 28590
rect 36990 28642 37042 28654
rect 42590 28642 42642 28654
rect 38546 28590 38558 28642
rect 38610 28590 38622 28642
rect 38994 28590 39006 28642
rect 39058 28590 39070 28642
rect 36990 28578 37042 28590
rect 42590 28578 42642 28590
rect 43934 28642 43986 28654
rect 43934 28578 43986 28590
rect 45054 28642 45106 28654
rect 45054 28578 45106 28590
rect 5966 28530 6018 28542
rect 5966 28466 6018 28478
rect 12910 28530 12962 28542
rect 12910 28466 12962 28478
rect 18398 28530 18450 28542
rect 18398 28466 18450 28478
rect 18510 28530 18562 28542
rect 18510 28466 18562 28478
rect 20638 28530 20690 28542
rect 27694 28530 27746 28542
rect 23538 28478 23550 28530
rect 23602 28478 23614 28530
rect 20638 28466 20690 28478
rect 27694 28466 27746 28478
rect 29486 28530 29538 28542
rect 29486 28466 29538 28478
rect 32734 28530 32786 28542
rect 32734 28466 32786 28478
rect 42926 28530 42978 28542
rect 42926 28466 42978 28478
rect 43150 28530 43202 28542
rect 43150 28466 43202 28478
rect 43374 28530 43426 28542
rect 43374 28466 43426 28478
rect 43486 28530 43538 28542
rect 43486 28466 43538 28478
rect 1710 28418 1762 28430
rect 18734 28418 18786 28430
rect 16370 28366 16382 28418
rect 16434 28366 16446 28418
rect 1710 28354 1762 28366
rect 18734 28354 18786 28366
rect 19182 28418 19234 28430
rect 19182 28354 19234 28366
rect 23214 28418 23266 28430
rect 42142 28418 42194 28430
rect 33730 28366 33742 28418
rect 33794 28366 33806 28418
rect 37314 28366 37326 28418
rect 37378 28366 37390 28418
rect 41570 28366 41582 28418
rect 41634 28366 41646 28418
rect 23214 28354 23266 28366
rect 42142 28354 42194 28366
rect 42814 28418 42866 28430
rect 42814 28354 42866 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 2046 28082 2098 28094
rect 2046 28018 2098 28030
rect 9886 28082 9938 28094
rect 9886 28018 9938 28030
rect 23214 28082 23266 28094
rect 23214 28018 23266 28030
rect 24670 28082 24722 28094
rect 24670 28018 24722 28030
rect 25566 28082 25618 28094
rect 25566 28018 25618 28030
rect 26014 28082 26066 28094
rect 31278 28082 31330 28094
rect 38894 28082 38946 28094
rect 27682 28030 27694 28082
rect 27746 28030 27758 28082
rect 35858 28030 35870 28082
rect 35922 28030 35934 28082
rect 36866 28030 36878 28082
rect 36930 28030 36942 28082
rect 44482 28030 44494 28082
rect 44546 28030 44558 28082
rect 26014 28018 26066 28030
rect 31278 28018 31330 28030
rect 38894 28018 38946 28030
rect 8318 27970 8370 27982
rect 18622 27970 18674 27982
rect 26126 27970 26178 27982
rect 17938 27918 17950 27970
rect 18002 27918 18014 27970
rect 22866 27918 22878 27970
rect 22930 27918 22942 27970
rect 8318 27906 8370 27918
rect 18622 27906 18674 27918
rect 26126 27906 26178 27918
rect 29598 27970 29650 27982
rect 54238 27970 54290 27982
rect 46386 27918 46398 27970
rect 46450 27918 46462 27970
rect 29598 27906 29650 27918
rect 54238 27906 54290 27918
rect 1710 27858 1762 27870
rect 1710 27794 1762 27806
rect 5630 27858 5682 27870
rect 9550 27858 9602 27870
rect 18846 27858 18898 27870
rect 6066 27806 6078 27858
rect 6130 27806 6142 27858
rect 18162 27806 18174 27858
rect 18226 27806 18238 27858
rect 5630 27794 5682 27806
rect 9550 27794 9602 27806
rect 18846 27794 18898 27806
rect 19406 27858 19458 27870
rect 19406 27794 19458 27806
rect 25230 27858 25282 27870
rect 25230 27794 25282 27806
rect 27134 27858 27186 27870
rect 30942 27858 30994 27870
rect 28466 27806 28478 27858
rect 28530 27806 28542 27858
rect 30034 27806 30046 27858
rect 30098 27806 30110 27858
rect 27134 27794 27186 27806
rect 30942 27794 30994 27806
rect 33182 27858 33234 27870
rect 36654 27858 36706 27870
rect 33618 27806 33630 27858
rect 33682 27806 33694 27858
rect 33182 27794 33234 27806
rect 36654 27794 36706 27806
rect 37214 27858 37266 27870
rect 37214 27794 37266 27806
rect 38558 27858 38610 27870
rect 38558 27794 38610 27806
rect 39006 27858 39058 27870
rect 39006 27794 39058 27806
rect 39230 27858 39282 27870
rect 39230 27794 39282 27806
rect 41358 27858 41410 27870
rect 49646 27858 49698 27870
rect 42018 27806 42030 27858
rect 42082 27806 42094 27858
rect 47282 27806 47294 27858
rect 47346 27806 47358 27858
rect 41358 27794 41410 27806
rect 49646 27794 49698 27806
rect 50430 27858 50482 27870
rect 50430 27794 50482 27806
rect 50878 27858 50930 27870
rect 50878 27794 50930 27806
rect 51102 27858 51154 27870
rect 53566 27858 53618 27870
rect 51986 27806 51998 27858
rect 52050 27806 52062 27858
rect 52882 27806 52894 27858
rect 52946 27806 52958 27858
rect 51102 27794 51154 27806
rect 53566 27794 53618 27806
rect 53902 27858 53954 27870
rect 53902 27794 53954 27806
rect 2494 27746 2546 27758
rect 2494 27682 2546 27694
rect 24222 27746 24274 27758
rect 24222 27682 24274 27694
rect 26910 27746 26962 27758
rect 31726 27746 31778 27758
rect 28130 27694 28142 27746
rect 28194 27694 28206 27746
rect 30482 27694 30494 27746
rect 30546 27694 30558 27746
rect 26910 27682 26962 27694
rect 31726 27682 31778 27694
rect 45390 27746 45442 27758
rect 47966 27746 48018 27758
rect 45826 27694 45838 27746
rect 45890 27694 45902 27746
rect 45390 27682 45442 27694
rect 47966 27682 48018 27694
rect 49422 27746 49474 27758
rect 49422 27682 49474 27694
rect 49870 27746 49922 27758
rect 49870 27682 49922 27694
rect 50990 27746 51042 27758
rect 50990 27682 51042 27694
rect 51438 27746 51490 27758
rect 53106 27694 53118 27746
rect 53170 27694 53182 27746
rect 51438 27682 51490 27694
rect 9102 27634 9154 27646
rect 9102 27570 9154 27582
rect 18734 27634 18786 27646
rect 18734 27570 18786 27582
rect 19182 27634 19234 27646
rect 19182 27570 19234 27582
rect 26014 27634 26066 27646
rect 26014 27570 26066 27582
rect 27358 27634 27410 27646
rect 27358 27570 27410 27582
rect 45054 27634 45106 27646
rect 45054 27570 45106 27582
rect 50318 27634 50370 27646
rect 50318 27570 50370 27582
rect 51662 27634 51714 27646
rect 51662 27570 51714 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 43262 27298 43314 27310
rect 43262 27234 43314 27246
rect 47406 27298 47458 27310
rect 47406 27234 47458 27246
rect 49086 27298 49138 27310
rect 49086 27234 49138 27246
rect 49758 27298 49810 27310
rect 49758 27234 49810 27246
rect 49982 27298 50034 27310
rect 49982 27234 50034 27246
rect 57934 27298 57986 27310
rect 57934 27234 57986 27246
rect 1934 27186 1986 27198
rect 1934 27122 1986 27134
rect 10334 27186 10386 27198
rect 10334 27122 10386 27134
rect 25678 27186 25730 27198
rect 25678 27122 25730 27134
rect 26686 27186 26738 27198
rect 26686 27122 26738 27134
rect 41022 27186 41074 27198
rect 41022 27122 41074 27134
rect 53118 27186 53170 27198
rect 53118 27122 53170 27134
rect 8878 27074 8930 27086
rect 18734 27074 18786 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 9650 27022 9662 27074
rect 9714 27022 9726 27074
rect 18386 27022 18398 27074
rect 18450 27022 18462 27074
rect 8878 27010 8930 27022
rect 18734 27010 18786 27022
rect 22766 27074 22818 27086
rect 46846 27074 46898 27086
rect 51774 27074 51826 27086
rect 33282 27022 33294 27074
rect 33346 27022 33358 27074
rect 34066 27022 34078 27074
rect 34130 27022 34142 27074
rect 37986 27022 37998 27074
rect 38050 27022 38062 27074
rect 41458 27022 41470 27074
rect 41522 27022 41534 27074
rect 45602 27022 45614 27074
rect 45666 27022 45678 27074
rect 49074 27022 49086 27074
rect 49138 27022 49150 27074
rect 49522 27022 49534 27074
rect 49586 27022 49598 27074
rect 22766 27010 22818 27022
rect 46846 27010 46898 27022
rect 51774 27010 51826 27022
rect 52558 27074 52610 27086
rect 55570 27022 55582 27074
rect 55634 27022 55646 27074
rect 52558 27010 52610 27022
rect 12462 26962 12514 26974
rect 9202 26910 9214 26962
rect 9266 26910 9278 26962
rect 9874 26910 9886 26962
rect 9938 26910 9950 26962
rect 12462 26898 12514 26910
rect 15038 26962 15090 26974
rect 15038 26898 15090 26910
rect 16046 26962 16098 26974
rect 16046 26898 16098 26910
rect 22654 26962 22706 26974
rect 22654 26898 22706 26910
rect 23326 26962 23378 26974
rect 23326 26898 23378 26910
rect 23438 26962 23490 26974
rect 23438 26898 23490 26910
rect 30830 26962 30882 26974
rect 30830 26898 30882 26910
rect 33518 26962 33570 26974
rect 33518 26898 33570 26910
rect 33854 26962 33906 26974
rect 33854 26898 33906 26910
rect 38222 26962 38274 26974
rect 43486 26962 43538 26974
rect 47070 26962 47122 26974
rect 38882 26910 38894 26962
rect 38946 26910 38958 26962
rect 45826 26910 45838 26962
rect 45890 26910 45902 26962
rect 38222 26898 38274 26910
rect 43486 26898 43538 26910
rect 47070 26898 47122 26910
rect 47294 26962 47346 26974
rect 47294 26898 47346 26910
rect 48750 26962 48802 26974
rect 48750 26898 48802 26910
rect 50094 26962 50146 26974
rect 50094 26898 50146 26910
rect 51438 26962 51490 26974
rect 51438 26898 51490 26910
rect 51662 26962 51714 26974
rect 51662 26898 51714 26910
rect 12126 26850 12178 26862
rect 12126 26786 12178 26798
rect 15262 26850 15314 26862
rect 15262 26786 15314 26798
rect 22878 26850 22930 26862
rect 22878 26786 22930 26798
rect 23662 26850 23714 26862
rect 23662 26786 23714 26798
rect 40686 26850 40738 26862
rect 40686 26786 40738 26798
rect 43374 26850 43426 26862
rect 43374 26786 43426 26798
rect 46174 26850 46226 26862
rect 46174 26786 46226 26798
rect 46286 26850 46338 26862
rect 46286 26786 46338 26798
rect 46398 26850 46450 26862
rect 46398 26786 46450 26798
rect 53006 26850 53058 26862
rect 53006 26786 53058 26798
rect 53230 26850 53282 26862
rect 53230 26786 53282 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 2046 26514 2098 26526
rect 2046 26450 2098 26462
rect 2718 26514 2770 26526
rect 36542 26514 36594 26526
rect 5058 26462 5070 26514
rect 5122 26462 5134 26514
rect 2718 26450 2770 26462
rect 36542 26450 36594 26462
rect 38558 26514 38610 26526
rect 38558 26450 38610 26462
rect 38782 26514 38834 26526
rect 38782 26450 38834 26462
rect 39566 26514 39618 26526
rect 39566 26450 39618 26462
rect 40238 26514 40290 26526
rect 40238 26450 40290 26462
rect 42142 26514 42194 26526
rect 42142 26450 42194 26462
rect 43374 26514 43426 26526
rect 43374 26450 43426 26462
rect 46510 26514 46562 26526
rect 46510 26450 46562 26462
rect 47070 26514 47122 26526
rect 47070 26450 47122 26462
rect 1710 26402 1762 26414
rect 1710 26338 1762 26350
rect 8206 26402 8258 26414
rect 8206 26338 8258 26350
rect 9662 26402 9714 26414
rect 9662 26338 9714 26350
rect 9998 26402 10050 26414
rect 9998 26338 10050 26350
rect 21198 26402 21250 26414
rect 21198 26338 21250 26350
rect 22542 26402 22594 26414
rect 22542 26338 22594 26350
rect 28366 26402 28418 26414
rect 36878 26402 36930 26414
rect 36194 26350 36206 26402
rect 36258 26350 36270 26402
rect 28366 26338 28418 26350
rect 36878 26338 36930 26350
rect 39678 26402 39730 26414
rect 39678 26338 39730 26350
rect 40350 26402 40402 26414
rect 40350 26338 40402 26350
rect 43038 26402 43090 26414
rect 43038 26338 43090 26350
rect 43150 26402 43202 26414
rect 43150 26338 43202 26350
rect 45838 26402 45890 26414
rect 45838 26338 45890 26350
rect 45950 26402 46002 26414
rect 45950 26338 46002 26350
rect 46286 26402 46338 26414
rect 46286 26338 46338 26350
rect 46622 26402 46674 26414
rect 46622 26338 46674 26350
rect 49758 26402 49810 26414
rect 49758 26338 49810 26350
rect 50318 26402 50370 26414
rect 50318 26338 50370 26350
rect 55022 26402 55074 26414
rect 55022 26338 55074 26350
rect 2382 26290 2434 26302
rect 2382 26226 2434 26238
rect 4398 26290 4450 26302
rect 5518 26290 5570 26302
rect 23774 26290 23826 26302
rect 4834 26238 4846 26290
rect 4898 26238 4910 26290
rect 5954 26238 5966 26290
rect 6018 26238 6030 26290
rect 10434 26238 10446 26290
rect 10498 26238 10510 26290
rect 11218 26238 11230 26290
rect 11282 26238 11294 26290
rect 11778 26238 11790 26290
rect 11842 26238 11854 26290
rect 14018 26238 14030 26290
rect 14082 26238 14094 26290
rect 20066 26238 20078 26290
rect 20130 26238 20142 26290
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 22978 26238 22990 26290
rect 23042 26238 23054 26290
rect 4398 26226 4450 26238
rect 5518 26226 5570 26238
rect 23774 26226 23826 26238
rect 24222 26290 24274 26302
rect 24222 26226 24274 26238
rect 24334 26290 24386 26302
rect 28254 26290 28306 26302
rect 25890 26238 25902 26290
rect 25954 26238 25966 26290
rect 26114 26238 26126 26290
rect 26178 26238 26190 26290
rect 24334 26226 24386 26238
rect 28254 26226 28306 26238
rect 39230 26290 39282 26302
rect 39230 26226 39282 26238
rect 40014 26290 40066 26302
rect 40014 26226 40066 26238
rect 43710 26290 43762 26302
rect 43710 26226 43762 26238
rect 48862 26290 48914 26302
rect 50206 26290 50258 26302
rect 49074 26238 49086 26290
rect 49138 26238 49150 26290
rect 48862 26226 48914 26238
rect 50206 26226 50258 26238
rect 50542 26290 50594 26302
rect 53006 26290 53058 26302
rect 54350 26290 54402 26302
rect 50754 26238 50766 26290
rect 50818 26238 50830 26290
rect 50978 26238 50990 26290
rect 51042 26238 51054 26290
rect 51986 26238 51998 26290
rect 52050 26238 52062 26290
rect 52322 26238 52334 26290
rect 52386 26238 52398 26290
rect 53666 26238 53678 26290
rect 53730 26238 53742 26290
rect 50542 26226 50594 26238
rect 53006 26226 53058 26238
rect 54350 26226 54402 26238
rect 54686 26290 54738 26302
rect 54686 26226 54738 26238
rect 3166 26178 3218 26190
rect 19630 26178 19682 26190
rect 23998 26178 24050 26190
rect 26910 26178 26962 26190
rect 10770 26126 10782 26178
rect 10834 26126 10846 26178
rect 20402 26126 20414 26178
rect 20466 26126 20478 26178
rect 22082 26126 22094 26178
rect 22146 26126 22158 26178
rect 23314 26126 23326 26178
rect 23378 26126 23390 26178
rect 26002 26126 26014 26178
rect 26066 26126 26078 26178
rect 3166 26114 3218 26126
rect 19630 26114 19682 26126
rect 23998 26114 24050 26126
rect 26910 26114 26962 26126
rect 27470 26178 27522 26190
rect 27470 26114 27522 26126
rect 29038 26178 29090 26190
rect 29038 26114 29090 26126
rect 31054 26178 31106 26190
rect 31054 26114 31106 26126
rect 38222 26178 38274 26190
rect 38222 26114 38274 26126
rect 38670 26178 38722 26190
rect 38670 26114 38722 26126
rect 42702 26178 42754 26190
rect 42702 26114 42754 26126
rect 46958 26178 47010 26190
rect 53554 26126 53566 26178
rect 53618 26126 53630 26178
rect 46958 26114 47010 26126
rect 8990 26066 9042 26078
rect 28366 26066 28418 26078
rect 15026 26014 15038 26066
rect 15090 26014 15102 26066
rect 25330 26014 25342 26066
rect 25394 26014 25406 26066
rect 8990 26002 9042 26014
rect 28366 26002 28418 26014
rect 36990 26066 37042 26078
rect 36990 26002 37042 26014
rect 39454 26066 39506 26078
rect 39454 26002 39506 26014
rect 45950 26066 46002 26078
rect 50754 26014 50766 26066
rect 50818 26014 50830 26066
rect 45950 26002 46002 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 22878 25730 22930 25742
rect 22530 25678 22542 25730
rect 22594 25678 22606 25730
rect 22878 25666 22930 25678
rect 29710 25730 29762 25742
rect 29710 25666 29762 25678
rect 52782 25730 52834 25742
rect 52782 25666 52834 25678
rect 57934 25730 57986 25742
rect 57934 25666 57986 25678
rect 2494 25618 2546 25630
rect 2494 25554 2546 25566
rect 5742 25618 5794 25630
rect 5742 25554 5794 25566
rect 15262 25618 15314 25630
rect 15262 25554 15314 25566
rect 20302 25618 20354 25630
rect 20302 25554 20354 25566
rect 20414 25618 20466 25630
rect 20414 25554 20466 25566
rect 21422 25618 21474 25630
rect 21422 25554 21474 25566
rect 23102 25618 23154 25630
rect 23102 25554 23154 25566
rect 23774 25618 23826 25630
rect 23774 25554 23826 25566
rect 24670 25618 24722 25630
rect 37886 25618 37938 25630
rect 30818 25566 30830 25618
rect 30882 25566 30894 25618
rect 35522 25566 35534 25618
rect 35586 25566 35598 25618
rect 24670 25554 24722 25566
rect 37886 25554 37938 25566
rect 42590 25618 42642 25630
rect 42590 25554 42642 25566
rect 43486 25618 43538 25630
rect 43486 25554 43538 25566
rect 47182 25618 47234 25630
rect 47182 25554 47234 25566
rect 51550 25618 51602 25630
rect 51550 25554 51602 25566
rect 52670 25618 52722 25630
rect 52670 25554 52722 25566
rect 5070 25506 5122 25518
rect 4162 25454 4174 25506
rect 4226 25454 4238 25506
rect 5070 25442 5122 25454
rect 6526 25506 6578 25518
rect 14030 25506 14082 25518
rect 17838 25506 17890 25518
rect 18734 25506 18786 25518
rect 25342 25506 25394 25518
rect 29486 25506 29538 25518
rect 8754 25454 8766 25506
rect 8818 25454 8830 25506
rect 9202 25454 9214 25506
rect 9266 25454 9278 25506
rect 11330 25454 11342 25506
rect 11394 25454 11406 25506
rect 14466 25454 14478 25506
rect 14530 25454 14542 25506
rect 18274 25454 18286 25506
rect 18338 25454 18350 25506
rect 20626 25454 20638 25506
rect 20690 25454 20702 25506
rect 27906 25454 27918 25506
rect 27970 25454 27982 25506
rect 6526 25442 6578 25454
rect 14030 25442 14082 25454
rect 17838 25442 17890 25454
rect 18734 25442 18786 25454
rect 25342 25442 25394 25454
rect 29486 25442 29538 25454
rect 29934 25506 29986 25518
rect 29934 25442 29986 25454
rect 30382 25506 30434 25518
rect 30382 25442 30434 25454
rect 31278 25506 31330 25518
rect 33742 25506 33794 25518
rect 31490 25454 31502 25506
rect 31554 25454 31566 25506
rect 32834 25454 32846 25506
rect 32898 25454 32910 25506
rect 33394 25454 33406 25506
rect 33458 25454 33470 25506
rect 31278 25442 31330 25454
rect 33742 25442 33794 25454
rect 34078 25506 34130 25518
rect 42366 25506 42418 25518
rect 35186 25454 35198 25506
rect 35250 25454 35262 25506
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 39554 25454 39566 25506
rect 39618 25454 39630 25506
rect 34078 25442 34130 25454
rect 42366 25442 42418 25454
rect 42702 25506 42754 25518
rect 42702 25442 42754 25454
rect 43038 25506 43090 25518
rect 43038 25442 43090 25454
rect 46286 25506 46338 25518
rect 50654 25506 50706 25518
rect 46498 25454 46510 25506
rect 46562 25454 46574 25506
rect 50866 25454 50878 25506
rect 50930 25454 50942 25506
rect 55570 25454 55582 25506
rect 55634 25454 55646 25506
rect 46286 25442 46338 25454
rect 50654 25442 50706 25454
rect 1710 25394 1762 25406
rect 1710 25330 1762 25342
rect 2046 25394 2098 25406
rect 2046 25330 2098 25342
rect 4398 25394 4450 25406
rect 4398 25330 4450 25342
rect 6190 25394 6242 25406
rect 6190 25330 6242 25342
rect 15374 25394 15426 25406
rect 15374 25330 15426 25342
rect 16046 25394 16098 25406
rect 16046 25330 16098 25342
rect 16606 25394 16658 25406
rect 16606 25330 16658 25342
rect 24782 25394 24834 25406
rect 24782 25330 24834 25342
rect 27582 25394 27634 25406
rect 32062 25394 32114 25406
rect 43374 25394 43426 25406
rect 28242 25342 28254 25394
rect 28306 25342 28318 25394
rect 40226 25342 40238 25394
rect 40290 25342 40302 25394
rect 27582 25330 27634 25342
rect 32062 25330 32114 25342
rect 43374 25330 43426 25342
rect 2942 25282 2994 25294
rect 17614 25282 17666 25294
rect 4722 25230 4734 25282
rect 4786 25230 4798 25282
rect 12450 25230 12462 25282
rect 12514 25230 12526 25282
rect 2942 25218 2994 25230
rect 17614 25218 17666 25230
rect 19406 25282 19458 25294
rect 19406 25218 19458 25230
rect 25006 25282 25058 25294
rect 25006 25218 25058 25230
rect 27246 25282 27298 25294
rect 27246 25218 27298 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 28590 25282 28642 25294
rect 28590 25218 28642 25230
rect 29038 25282 29090 25294
rect 29038 25218 29090 25230
rect 34302 25282 34354 25294
rect 37326 25282 37378 25294
rect 34626 25230 34638 25282
rect 34690 25230 34702 25282
rect 34302 25218 34354 25230
rect 37326 25218 37378 25230
rect 43598 25282 43650 25294
rect 43598 25218 43650 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 20862 24946 20914 24958
rect 20862 24882 20914 24894
rect 25790 24946 25842 24958
rect 25790 24882 25842 24894
rect 34190 24946 34242 24958
rect 34190 24882 34242 24894
rect 42142 24946 42194 24958
rect 42142 24882 42194 24894
rect 48862 24946 48914 24958
rect 48862 24882 48914 24894
rect 53006 24946 53058 24958
rect 53006 24882 53058 24894
rect 23662 24834 23714 24846
rect 19282 24782 19294 24834
rect 19346 24782 19358 24834
rect 17390 24722 17442 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 5058 24670 5070 24722
rect 5122 24670 5134 24722
rect 5506 24670 5518 24722
rect 5570 24670 5582 24722
rect 7746 24670 7758 24722
rect 7810 24670 7822 24722
rect 14130 24670 14142 24722
rect 14194 24670 14206 24722
rect 15250 24670 15262 24722
rect 15314 24670 15326 24722
rect 16370 24670 16382 24722
rect 16434 24670 16446 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 17390 24658 17442 24670
rect 12686 24610 12738 24622
rect 12686 24546 12738 24558
rect 13918 24610 13970 24622
rect 13918 24546 13970 24558
rect 18510 24610 18562 24622
rect 18510 24546 18562 24558
rect 19070 24610 19122 24622
rect 19070 24546 19122 24558
rect 1934 24498 1986 24510
rect 8754 24446 8766 24498
rect 8818 24446 8830 24498
rect 16258 24446 16270 24498
rect 16322 24446 16334 24498
rect 18722 24446 18734 24498
rect 18786 24495 18798 24498
rect 19297 24495 19343 24782
rect 23662 24770 23714 24782
rect 29822 24834 29874 24846
rect 34414 24834 34466 24846
rect 33618 24782 33630 24834
rect 33682 24782 33694 24834
rect 29822 24770 29874 24782
rect 34414 24770 34466 24782
rect 35646 24834 35698 24846
rect 49646 24834 49698 24846
rect 41794 24782 41806 24834
rect 41858 24782 41870 24834
rect 43362 24782 43374 24834
rect 43426 24782 43438 24834
rect 35646 24770 35698 24782
rect 49646 24770 49698 24782
rect 19854 24722 19906 24734
rect 26910 24722 26962 24734
rect 23090 24670 23102 24722
rect 23154 24670 23166 24722
rect 26002 24670 26014 24722
rect 26066 24670 26078 24722
rect 19854 24658 19906 24670
rect 26910 24658 26962 24670
rect 28142 24722 28194 24734
rect 30718 24722 30770 24734
rect 28466 24670 28478 24722
rect 28530 24670 28542 24722
rect 28142 24658 28194 24670
rect 30718 24658 30770 24670
rect 30830 24722 30882 24734
rect 30830 24658 30882 24670
rect 31166 24722 31218 24734
rect 31166 24658 31218 24670
rect 32062 24722 32114 24734
rect 32062 24658 32114 24670
rect 33294 24722 33346 24734
rect 33294 24658 33346 24670
rect 33854 24722 33906 24734
rect 33854 24658 33906 24670
rect 35086 24722 35138 24734
rect 47070 24722 47122 24734
rect 35410 24670 35422 24722
rect 35474 24670 35486 24722
rect 43138 24670 43150 24722
rect 43202 24670 43214 24722
rect 44706 24670 44718 24722
rect 44770 24670 44782 24722
rect 46274 24670 46286 24722
rect 46338 24670 46350 24722
rect 35086 24658 35138 24670
rect 47070 24658 47122 24670
rect 48750 24722 48802 24734
rect 48750 24658 48802 24670
rect 48974 24722 49026 24734
rect 48974 24658 49026 24670
rect 49422 24722 49474 24734
rect 49422 24658 49474 24670
rect 52894 24722 52946 24734
rect 52894 24658 52946 24670
rect 53230 24722 53282 24734
rect 53890 24670 53902 24722
rect 53954 24670 53966 24722
rect 53230 24658 53282 24670
rect 19518 24610 19570 24622
rect 19518 24546 19570 24558
rect 20414 24610 20466 24622
rect 20414 24546 20466 24558
rect 22878 24610 22930 24622
rect 22878 24546 22930 24558
rect 25342 24610 25394 24622
rect 25342 24546 25394 24558
rect 25678 24610 25730 24622
rect 31054 24610 31106 24622
rect 26450 24558 26462 24610
rect 26514 24558 26526 24610
rect 28690 24558 28702 24610
rect 28754 24558 28766 24610
rect 25678 24546 25730 24558
rect 31054 24546 31106 24558
rect 31726 24610 31778 24622
rect 31726 24546 31778 24558
rect 34526 24610 34578 24622
rect 34526 24546 34578 24558
rect 34862 24610 34914 24622
rect 34862 24546 34914 24558
rect 36430 24610 36482 24622
rect 36430 24546 36482 24558
rect 36990 24610 37042 24622
rect 44370 24558 44382 24610
rect 44434 24558 44446 24610
rect 36990 24546 37042 24558
rect 18786 24449 19343 24495
rect 23326 24498 23378 24510
rect 18786 24446 18798 24449
rect 1934 24434 1986 24446
rect 23326 24434 23378 24446
rect 23550 24498 23602 24510
rect 29934 24498 29986 24510
rect 35758 24498 35810 24510
rect 49758 24498 49810 24510
rect 28466 24446 28478 24498
rect 28530 24446 28542 24498
rect 34626 24446 34638 24498
rect 34690 24495 34702 24498
rect 34962 24495 34974 24498
rect 34690 24449 34974 24495
rect 34690 24446 34702 24449
rect 34962 24446 34974 24449
rect 35026 24446 35038 24498
rect 36306 24446 36318 24498
rect 36370 24495 36382 24498
rect 36978 24495 36990 24498
rect 36370 24449 36990 24495
rect 36370 24446 36382 24449
rect 36978 24446 36990 24449
rect 37042 24446 37054 24498
rect 55346 24446 55358 24498
rect 55410 24446 55422 24498
rect 23550 24434 23602 24446
rect 29934 24434 29986 24446
rect 35758 24434 35810 24446
rect 49758 24434 49810 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 19518 24162 19570 24174
rect 18274 24110 18286 24162
rect 18338 24110 18350 24162
rect 19518 24098 19570 24110
rect 35646 24162 35698 24174
rect 35646 24098 35698 24110
rect 43150 24162 43202 24174
rect 43150 24098 43202 24110
rect 43486 24162 43538 24174
rect 57934 24162 57986 24174
rect 46834 24110 46846 24162
rect 46898 24110 46910 24162
rect 53666 24110 53678 24162
rect 53730 24110 53742 24162
rect 43486 24098 43538 24110
rect 57934 24098 57986 24110
rect 1934 24050 1986 24062
rect 10446 24050 10498 24062
rect 15934 24050 15986 24062
rect 30046 24050 30098 24062
rect 42478 24050 42530 24062
rect 9538 23998 9550 24050
rect 9602 23998 9614 24050
rect 10882 23998 10894 24050
rect 10946 23998 10958 24050
rect 11890 23998 11902 24050
rect 11954 23998 11966 24050
rect 16258 23998 16270 24050
rect 16322 23998 16334 24050
rect 25218 23998 25230 24050
rect 25282 23998 25294 24050
rect 28354 23998 28366 24050
rect 28418 23998 28430 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 45602 23998 45614 24050
rect 45666 23998 45678 24050
rect 46946 23998 46958 24050
rect 47010 23998 47022 24050
rect 48178 23998 48190 24050
rect 48242 23998 48254 24050
rect 49298 23998 49310 24050
rect 49362 23998 49374 24050
rect 53330 23998 53342 24050
rect 53394 23998 53406 24050
rect 1934 23986 1986 23998
rect 10446 23986 10498 23998
rect 15934 23986 15986 23998
rect 30046 23986 30098 23998
rect 42478 23986 42530 23998
rect 5966 23938 6018 23950
rect 14366 23938 14418 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 11218 23886 11230 23938
rect 11282 23886 11294 23938
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 5966 23874 6018 23886
rect 14366 23874 14418 23886
rect 14926 23938 14978 23950
rect 14926 23874 14978 23886
rect 15374 23938 15426 23950
rect 19294 23938 19346 23950
rect 16482 23886 16494 23938
rect 16546 23886 16558 23938
rect 18610 23886 18622 23938
rect 18674 23886 18686 23938
rect 15374 23874 15426 23886
rect 19294 23874 19346 23886
rect 22990 23938 23042 23950
rect 30494 23938 30546 23950
rect 35758 23938 35810 23950
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 26114 23886 26126 23938
rect 26178 23886 26190 23938
rect 27122 23886 27134 23938
rect 27186 23886 27198 23938
rect 28130 23886 28142 23938
rect 28194 23886 28206 23938
rect 30930 23886 30942 23938
rect 30994 23886 31006 23938
rect 31714 23886 31726 23938
rect 31778 23886 31790 23938
rect 33394 23886 33406 23938
rect 33458 23886 33470 23938
rect 34738 23886 34750 23938
rect 34802 23886 34814 23938
rect 22990 23874 23042 23886
rect 30494 23874 30546 23886
rect 35758 23874 35810 23886
rect 36206 23938 36258 23950
rect 45166 23938 45218 23950
rect 48862 23938 48914 23950
rect 37090 23886 37102 23938
rect 37154 23886 37166 23938
rect 38770 23886 38782 23938
rect 38834 23886 38846 23938
rect 40786 23886 40798 23938
rect 40850 23886 40862 23938
rect 46050 23886 46062 23938
rect 46114 23886 46126 23938
rect 46722 23886 46734 23938
rect 46786 23886 46798 23938
rect 47954 23886 47966 23938
rect 48018 23886 48030 23938
rect 49746 23886 49758 23938
rect 49810 23886 49822 23938
rect 52882 23886 52894 23938
rect 52946 23886 52958 23938
rect 53442 23886 53454 23938
rect 53506 23886 53518 23938
rect 54674 23886 54686 23938
rect 54738 23886 54750 23938
rect 55570 23886 55582 23938
rect 55634 23886 55646 23938
rect 36206 23874 36258 23886
rect 45166 23874 45218 23886
rect 48862 23874 48914 23886
rect 5630 23826 5682 23838
rect 5630 23762 5682 23774
rect 22878 23826 22930 23838
rect 25006 23826 25058 23838
rect 23762 23774 23774 23826
rect 23826 23774 23838 23826
rect 22878 23762 22930 23774
rect 25006 23762 25058 23774
rect 25566 23826 25618 23838
rect 30270 23826 30322 23838
rect 44830 23826 44882 23838
rect 27570 23774 27582 23826
rect 27634 23774 27646 23826
rect 28018 23774 28030 23826
rect 28082 23774 28094 23826
rect 31826 23774 31838 23826
rect 31890 23774 31902 23826
rect 37874 23774 37886 23826
rect 37938 23774 37950 23826
rect 40338 23774 40350 23826
rect 40402 23774 40414 23826
rect 25566 23762 25618 23774
rect 30270 23762 30322 23774
rect 44830 23762 44882 23774
rect 50206 23826 50258 23838
rect 50206 23762 50258 23774
rect 54462 23826 54514 23838
rect 54462 23762 54514 23774
rect 9102 23714 9154 23726
rect 9102 23650 9154 23662
rect 12350 23714 12402 23726
rect 12350 23650 12402 23662
rect 12798 23714 12850 23726
rect 12798 23650 12850 23662
rect 15038 23714 15090 23726
rect 20526 23714 20578 23726
rect 19842 23662 19854 23714
rect 19906 23662 19918 23714
rect 15038 23650 15090 23662
rect 20526 23650 20578 23662
rect 21534 23714 21586 23726
rect 21534 23650 21586 23662
rect 21982 23714 22034 23726
rect 21982 23650 22034 23662
rect 22654 23714 22706 23726
rect 22654 23650 22706 23662
rect 23102 23714 23154 23726
rect 23102 23650 23154 23662
rect 24334 23714 24386 23726
rect 24334 23650 24386 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 29486 23714 29538 23726
rect 29486 23650 29538 23662
rect 30606 23714 30658 23726
rect 30606 23650 30658 23662
rect 30718 23714 30770 23726
rect 30718 23650 30770 23662
rect 35646 23714 35698 23726
rect 35646 23650 35698 23662
rect 41246 23714 41298 23726
rect 41246 23650 41298 23662
rect 42030 23714 42082 23726
rect 42030 23650 42082 23662
rect 42590 23714 42642 23726
rect 42590 23650 42642 23662
rect 43374 23714 43426 23726
rect 43374 23650 43426 23662
rect 44270 23714 44322 23726
rect 44270 23650 44322 23662
rect 44942 23714 44994 23726
rect 44942 23650 44994 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 12462 23378 12514 23390
rect 12462 23314 12514 23326
rect 17390 23378 17442 23390
rect 17390 23314 17442 23326
rect 18510 23378 18562 23390
rect 21422 23378 21474 23390
rect 20962 23326 20974 23378
rect 21026 23326 21038 23378
rect 18510 23314 18562 23326
rect 21422 23314 21474 23326
rect 24558 23378 24610 23390
rect 24558 23314 24610 23326
rect 26910 23378 26962 23390
rect 26910 23314 26962 23326
rect 34414 23378 34466 23390
rect 34414 23314 34466 23326
rect 35422 23378 35474 23390
rect 35422 23314 35474 23326
rect 36206 23378 36258 23390
rect 36206 23314 36258 23326
rect 36766 23378 36818 23390
rect 36766 23314 36818 23326
rect 36878 23378 36930 23390
rect 36878 23314 36930 23326
rect 38558 23378 38610 23390
rect 38558 23314 38610 23326
rect 44382 23378 44434 23390
rect 44382 23314 44434 23326
rect 49534 23378 49586 23390
rect 49534 23314 49586 23326
rect 51438 23378 51490 23390
rect 52670 23378 52722 23390
rect 52210 23326 52222 23378
rect 52274 23326 52286 23378
rect 51438 23314 51490 23326
rect 52670 23314 52722 23326
rect 53006 23378 53058 23390
rect 53006 23314 53058 23326
rect 12574 23266 12626 23278
rect 25566 23266 25618 23278
rect 8978 23214 8990 23266
rect 9042 23214 9054 23266
rect 12002 23214 12014 23266
rect 12066 23214 12078 23266
rect 13682 23214 13694 23266
rect 13746 23214 13758 23266
rect 12574 23202 12626 23214
rect 25566 23202 25618 23214
rect 32510 23266 32562 23278
rect 42366 23266 42418 23278
rect 37650 23214 37662 23266
rect 37714 23214 37726 23266
rect 37986 23214 37998 23266
rect 38050 23214 38062 23266
rect 41010 23214 41022 23266
rect 41074 23214 41086 23266
rect 41794 23214 41806 23266
rect 41858 23214 41870 23266
rect 32510 23202 32562 23214
rect 42366 23202 42418 23214
rect 44830 23266 44882 23278
rect 44830 23202 44882 23214
rect 49198 23266 49250 23278
rect 49198 23202 49250 23214
rect 49310 23266 49362 23278
rect 49310 23202 49362 23214
rect 51102 23266 51154 23278
rect 51102 23202 51154 23214
rect 51214 23266 51266 23278
rect 51214 23202 51266 23214
rect 51662 23266 51714 23278
rect 51662 23202 51714 23214
rect 54462 23266 54514 23278
rect 54462 23202 54514 23214
rect 8318 23154 8370 23166
rect 10558 23154 10610 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 7858 23102 7870 23154
rect 7922 23102 7934 23154
rect 8754 23102 8766 23154
rect 8818 23102 8830 23154
rect 10098 23102 10110 23154
rect 10162 23102 10174 23154
rect 8318 23090 8370 23102
rect 10558 23090 10610 23102
rect 11454 23154 11506 23166
rect 19854 23154 19906 23166
rect 13346 23102 13358 23154
rect 13410 23102 13422 23154
rect 16258 23102 16270 23154
rect 16322 23102 16334 23154
rect 16706 23102 16718 23154
rect 16770 23102 16782 23154
rect 11454 23090 11506 23102
rect 19854 23090 19906 23102
rect 20302 23154 20354 23166
rect 20302 23090 20354 23102
rect 20638 23154 20690 23166
rect 26350 23154 26402 23166
rect 27022 23154 27074 23166
rect 22754 23102 22766 23154
rect 22818 23102 22830 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 20638 23090 20690 23102
rect 26350 23090 26402 23102
rect 27022 23090 27074 23102
rect 27470 23154 27522 23166
rect 27470 23090 27522 23102
rect 27694 23154 27746 23166
rect 27694 23090 27746 23102
rect 28366 23154 28418 23166
rect 29934 23154 29986 23166
rect 30942 23154 30994 23166
rect 28578 23102 28590 23154
rect 28642 23102 28654 23154
rect 29586 23102 29598 23154
rect 29650 23102 29662 23154
rect 30370 23102 30382 23154
rect 30434 23102 30446 23154
rect 28366 23090 28418 23102
rect 29934 23090 29986 23102
rect 30942 23090 30994 23102
rect 31390 23154 31442 23166
rect 31390 23090 31442 23102
rect 31502 23154 31554 23166
rect 31502 23090 31554 23102
rect 31614 23154 31666 23166
rect 31614 23090 31666 23102
rect 34190 23154 34242 23166
rect 34190 23090 34242 23102
rect 34302 23154 34354 23166
rect 34302 23090 34354 23102
rect 34526 23154 34578 23166
rect 40126 23154 40178 23166
rect 42702 23154 42754 23166
rect 34738 23102 34750 23154
rect 34802 23102 34814 23154
rect 40898 23102 40910 23154
rect 40962 23102 40974 23154
rect 34526 23090 34578 23102
rect 40126 23090 40178 23102
rect 42702 23090 42754 23102
rect 44046 23154 44098 23166
rect 44046 23090 44098 23102
rect 44158 23154 44210 23166
rect 44158 23090 44210 23102
rect 44494 23154 44546 23166
rect 51886 23154 51938 23166
rect 45378 23102 45390 23154
rect 45442 23102 45454 23154
rect 44494 23090 44546 23102
rect 51886 23090 51938 23102
rect 52894 23154 52946 23166
rect 52894 23090 52946 23102
rect 53118 23154 53170 23166
rect 53778 23102 53790 23154
rect 53842 23102 53854 23154
rect 53118 23090 53170 23102
rect 17950 23042 18002 23054
rect 7970 22990 7982 23042
rect 8034 22990 8046 23042
rect 9762 22990 9774 23042
rect 9826 22990 9838 23042
rect 10994 22990 11006 23042
rect 11058 22990 11070 23042
rect 14578 22990 14590 23042
rect 14642 22990 14654 23042
rect 17950 22978 18002 22990
rect 19070 23042 19122 23054
rect 19070 22978 19122 22990
rect 19518 23042 19570 23054
rect 19518 22978 19570 22990
rect 21982 23042 22034 23054
rect 21982 22978 22034 22990
rect 22430 23042 22482 23054
rect 26126 23042 26178 23054
rect 22754 23039 22766 23042
rect 22430 22978 22482 22990
rect 22545 22993 22766 23039
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 11678 22930 11730 22942
rect 21858 22878 21870 22930
rect 21922 22927 21934 22930
rect 22545 22927 22591 22993
rect 22754 22990 22766 22993
rect 22818 22990 22830 23042
rect 23874 22990 23886 23042
rect 23938 22990 23950 23042
rect 25666 22990 25678 23042
rect 25730 22990 25742 23042
rect 26126 22978 26178 22990
rect 32174 23042 32226 23054
rect 32174 22978 32226 22990
rect 33742 23042 33794 23054
rect 33742 22978 33794 22990
rect 39006 23042 39058 23054
rect 39006 22978 39058 22990
rect 42142 23042 42194 23054
rect 42142 22978 42194 22990
rect 43150 23042 43202 23054
rect 47406 23042 47458 23054
rect 45602 22990 45614 23042
rect 45666 22990 45678 23042
rect 54002 22990 54014 23042
rect 54066 22990 54078 23042
rect 43150 22978 43202 22990
rect 47406 22978 47458 22990
rect 21922 22881 22591 22927
rect 25342 22930 25394 22942
rect 36654 22930 36706 22942
rect 21922 22878 21934 22881
rect 28018 22878 28030 22930
rect 28082 22878 28094 22930
rect 30034 22878 30046 22930
rect 30098 22878 30110 22930
rect 11678 22866 11730 22878
rect 25342 22866 25394 22878
rect 36654 22866 36706 22878
rect 38222 22930 38274 22942
rect 38222 22866 38274 22878
rect 39230 22930 39282 22942
rect 39230 22866 39282 22878
rect 39454 22930 39506 22942
rect 39454 22866 39506 22878
rect 39678 22930 39730 22942
rect 39678 22866 39730 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 37774 22594 37826 22606
rect 16482 22542 16494 22594
rect 16546 22542 16558 22594
rect 31266 22542 31278 22594
rect 31330 22542 31342 22594
rect 37774 22530 37826 22542
rect 39230 22594 39282 22606
rect 50766 22594 50818 22606
rect 47954 22542 47966 22594
rect 48018 22542 48030 22594
rect 39230 22530 39282 22542
rect 50766 22530 50818 22542
rect 1934 22482 1986 22494
rect 10894 22482 10946 22494
rect 27806 22482 27858 22494
rect 32622 22482 32674 22494
rect 8866 22430 8878 22482
rect 8930 22430 8942 22482
rect 16034 22430 16046 22482
rect 16098 22430 16110 22482
rect 20066 22430 20078 22482
rect 20130 22430 20142 22482
rect 30034 22430 30046 22482
rect 30098 22430 30110 22482
rect 31042 22430 31054 22482
rect 31106 22430 31118 22482
rect 1934 22418 1986 22430
rect 10894 22418 10946 22430
rect 27806 22418 27858 22430
rect 32622 22418 32674 22430
rect 36430 22482 36482 22494
rect 39006 22482 39058 22494
rect 54350 22482 54402 22494
rect 38098 22430 38110 22482
rect 38162 22430 38174 22482
rect 40002 22430 40014 22482
rect 40066 22430 40078 22482
rect 45378 22430 45390 22482
rect 45442 22430 45454 22482
rect 47282 22430 47294 22482
rect 47346 22430 47358 22482
rect 53778 22430 53790 22482
rect 53842 22430 53854 22482
rect 36430 22418 36482 22430
rect 39006 22418 39058 22430
rect 54350 22418 54402 22430
rect 9326 22370 9378 22382
rect 11230 22370 11282 22382
rect 4162 22318 4174 22370
rect 4226 22318 4238 22370
rect 9650 22318 9662 22370
rect 9714 22318 9726 22370
rect 9326 22306 9378 22318
rect 11230 22306 11282 22318
rect 11342 22370 11394 22382
rect 11342 22306 11394 22318
rect 11566 22370 11618 22382
rect 14254 22370 14306 22382
rect 13794 22318 13806 22370
rect 13858 22318 13870 22370
rect 11566 22306 11618 22318
rect 14254 22306 14306 22318
rect 14590 22370 14642 22382
rect 34974 22370 35026 22382
rect 15362 22318 15374 22370
rect 15426 22318 15438 22370
rect 16370 22318 16382 22370
rect 16434 22318 16446 22370
rect 17154 22318 17166 22370
rect 17218 22318 17230 22370
rect 19282 22318 19294 22370
rect 19346 22318 19358 22370
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 23650 22318 23662 22370
rect 23714 22318 23726 22370
rect 24770 22318 24782 22370
rect 24834 22318 24846 22370
rect 27458 22318 27470 22370
rect 27522 22318 27534 22370
rect 28242 22318 28254 22370
rect 28306 22318 28318 22370
rect 30258 22318 30270 22370
rect 30322 22318 30334 22370
rect 31378 22318 31390 22370
rect 31442 22318 31454 22370
rect 33058 22318 33070 22370
rect 33122 22318 33134 22370
rect 33954 22318 33966 22370
rect 34018 22318 34030 22370
rect 14590 22306 14642 22318
rect 34974 22306 35026 22318
rect 35310 22370 35362 22382
rect 35310 22306 35362 22318
rect 39454 22370 39506 22382
rect 40126 22370 40178 22382
rect 39778 22318 39790 22370
rect 39842 22318 39854 22370
rect 39454 22306 39506 22318
rect 40126 22306 40178 22318
rect 41358 22370 41410 22382
rect 41358 22306 41410 22318
rect 41582 22370 41634 22382
rect 41582 22306 41634 22318
rect 42030 22370 42082 22382
rect 42030 22306 42082 22318
rect 43710 22370 43762 22382
rect 43710 22306 43762 22318
rect 43822 22370 43874 22382
rect 50430 22370 50482 22382
rect 44706 22318 44718 22370
rect 44770 22318 44782 22370
rect 45490 22318 45502 22370
rect 45554 22318 45566 22370
rect 47506 22318 47518 22370
rect 47570 22318 47582 22370
rect 50194 22318 50206 22370
rect 50258 22318 50270 22370
rect 43822 22306 43874 22318
rect 50430 22306 50482 22318
rect 50654 22370 50706 22382
rect 53890 22318 53902 22370
rect 53954 22318 53966 22370
rect 50654 22306 50706 22318
rect 15150 22258 15202 22270
rect 18174 22258 18226 22270
rect 9762 22206 9774 22258
rect 9826 22206 9838 22258
rect 10210 22206 10222 22258
rect 10274 22206 10286 22258
rect 12114 22206 12126 22258
rect 12178 22206 12190 22258
rect 17266 22206 17278 22258
rect 17330 22206 17342 22258
rect 15150 22194 15202 22206
rect 18174 22194 18226 22206
rect 18286 22258 18338 22270
rect 32846 22258 32898 22270
rect 34526 22258 34578 22270
rect 20514 22206 20526 22258
rect 20578 22206 20590 22258
rect 21970 22206 21982 22258
rect 22034 22206 22046 22258
rect 25442 22206 25454 22258
rect 25506 22206 25518 22258
rect 26114 22206 26126 22258
rect 26178 22206 26190 22258
rect 27122 22206 27134 22258
rect 27186 22206 27198 22258
rect 27794 22206 27806 22258
rect 27858 22206 27870 22258
rect 34290 22206 34302 22258
rect 34354 22206 34366 22258
rect 18286 22194 18338 22206
rect 32846 22194 32898 22206
rect 34526 22194 34578 22206
rect 35534 22258 35586 22270
rect 35534 22194 35586 22206
rect 37998 22258 38050 22270
rect 37998 22194 38050 22206
rect 41806 22258 41858 22270
rect 41806 22194 41858 22206
rect 42142 22258 42194 22270
rect 53566 22258 53618 22270
rect 46162 22206 46174 22258
rect 46226 22206 46238 22258
rect 42142 22194 42194 22206
rect 53566 22194 53618 22206
rect 54238 22258 54290 22270
rect 54238 22194 54290 22206
rect 54462 22258 54514 22270
rect 54462 22194 54514 22206
rect 8430 22146 8482 22158
rect 8430 22082 8482 22094
rect 12910 22146 12962 22158
rect 18510 22146 18562 22158
rect 25790 22146 25842 22158
rect 17490 22094 17502 22146
rect 17554 22094 17566 22146
rect 25218 22094 25230 22146
rect 25282 22094 25294 22146
rect 12910 22082 12962 22094
rect 18510 22082 18562 22094
rect 25790 22082 25842 22094
rect 29374 22146 29426 22158
rect 29374 22082 29426 22094
rect 35422 22146 35474 22158
rect 35422 22082 35474 22094
rect 39902 22146 39954 22158
rect 39902 22082 39954 22094
rect 43038 22146 43090 22158
rect 43934 22146 43986 22158
rect 43362 22094 43374 22146
rect 43426 22094 43438 22146
rect 43038 22082 43090 22094
rect 43934 22082 43986 22094
rect 44158 22146 44210 22158
rect 44158 22082 44210 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 10782 21810 10834 21822
rect 6290 21758 6302 21810
rect 6354 21758 6366 21810
rect 10782 21746 10834 21758
rect 16046 21810 16098 21822
rect 16046 21746 16098 21758
rect 17390 21810 17442 21822
rect 17390 21746 17442 21758
rect 19294 21810 19346 21822
rect 19294 21746 19346 21758
rect 21758 21810 21810 21822
rect 21758 21746 21810 21758
rect 21982 21810 22034 21822
rect 21982 21746 22034 21758
rect 22878 21810 22930 21822
rect 22878 21746 22930 21758
rect 22990 21810 23042 21822
rect 27470 21810 27522 21822
rect 25330 21758 25342 21810
rect 25394 21758 25406 21810
rect 22990 21746 23042 21758
rect 27470 21746 27522 21758
rect 27694 21810 27746 21822
rect 27694 21746 27746 21758
rect 32622 21810 32674 21822
rect 32622 21746 32674 21758
rect 33406 21810 33458 21822
rect 33406 21746 33458 21758
rect 34974 21810 35026 21822
rect 44046 21810 44098 21822
rect 42802 21758 42814 21810
rect 42866 21758 42878 21810
rect 34974 21746 35026 21758
rect 44046 21746 44098 21758
rect 47518 21810 47570 21822
rect 47518 21746 47570 21758
rect 47630 21810 47682 21822
rect 47630 21746 47682 21758
rect 47742 21810 47794 21822
rect 47742 21746 47794 21758
rect 21646 21698 21698 21710
rect 6962 21646 6974 21698
rect 7026 21646 7038 21698
rect 16818 21646 16830 21698
rect 16882 21646 16894 21698
rect 20738 21646 20750 21698
rect 20802 21646 20814 21698
rect 21646 21634 21698 21646
rect 22206 21698 22258 21710
rect 22206 21634 22258 21646
rect 22318 21698 22370 21710
rect 27358 21698 27410 21710
rect 26674 21646 26686 21698
rect 26738 21646 26750 21698
rect 22318 21634 22370 21646
rect 27358 21634 27410 21646
rect 29150 21698 29202 21710
rect 29150 21634 29202 21646
rect 32398 21698 32450 21710
rect 34750 21698 34802 21710
rect 33058 21646 33070 21698
rect 33122 21646 33134 21698
rect 32398 21634 32450 21646
rect 34750 21634 34802 21646
rect 36878 21698 36930 21710
rect 41022 21698 41074 21710
rect 44158 21698 44210 21710
rect 37538 21646 37550 21698
rect 37602 21646 37614 21698
rect 42242 21646 42254 21698
rect 42306 21646 42318 21698
rect 36878 21634 36930 21646
rect 41022 21634 41074 21646
rect 44158 21634 44210 21646
rect 44830 21698 44882 21710
rect 44830 21634 44882 21646
rect 46734 21698 46786 21710
rect 54014 21698 54066 21710
rect 49410 21646 49422 21698
rect 49474 21646 49486 21698
rect 46734 21634 46786 21646
rect 54014 21634 54066 21646
rect 54574 21698 54626 21710
rect 54574 21634 54626 21646
rect 5966 21586 6018 21598
rect 15150 21586 15202 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 6738 21534 6750 21586
rect 6802 21534 6814 21586
rect 11554 21534 11566 21586
rect 11618 21534 11630 21586
rect 14130 21534 14142 21586
rect 14194 21534 14206 21586
rect 5966 21522 6018 21534
rect 15150 21522 15202 21534
rect 16494 21586 16546 21598
rect 16494 21522 16546 21534
rect 17950 21586 18002 21598
rect 23102 21586 23154 21598
rect 24110 21586 24162 21598
rect 19618 21534 19630 21586
rect 19682 21534 19694 21586
rect 22642 21534 22654 21586
rect 22706 21534 22718 21586
rect 23314 21534 23326 21586
rect 23378 21534 23390 21586
rect 17950 21522 18002 21534
rect 23102 21522 23154 21534
rect 24110 21522 24162 21534
rect 24334 21586 24386 21598
rect 24334 21522 24386 21534
rect 24670 21586 24722 21598
rect 28366 21586 28418 21598
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 26114 21534 26126 21586
rect 26178 21534 26190 21586
rect 24670 21522 24722 21534
rect 28366 21522 28418 21534
rect 28814 21586 28866 21598
rect 30830 21586 30882 21598
rect 32286 21586 32338 21598
rect 34638 21586 34690 21598
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 30146 21534 30158 21586
rect 30210 21534 30222 21586
rect 31042 21534 31054 21586
rect 31106 21534 31118 21586
rect 34178 21534 34190 21586
rect 34242 21534 34254 21586
rect 28814 21522 28866 21534
rect 30830 21522 30882 21534
rect 32286 21522 32338 21534
rect 34638 21522 34690 21534
rect 35982 21586 36034 21598
rect 38110 21586 38162 21598
rect 43486 21586 43538 21598
rect 36194 21534 36206 21586
rect 36258 21534 36270 21586
rect 37314 21534 37326 21586
rect 37378 21534 37390 21586
rect 42130 21534 42142 21586
rect 42194 21534 42206 21586
rect 42802 21534 42814 21586
rect 42866 21534 42878 21586
rect 35982 21522 36034 21534
rect 38110 21522 38162 21534
rect 43486 21522 43538 21534
rect 43710 21586 43762 21598
rect 43710 21522 43762 21534
rect 44382 21586 44434 21598
rect 44382 21522 44434 21534
rect 46846 21586 46898 21598
rect 46846 21522 46898 21534
rect 47070 21586 47122 21598
rect 49746 21534 49758 21586
rect 49810 21534 49822 21586
rect 50866 21534 50878 21586
rect 50930 21534 50942 21586
rect 53106 21534 53118 21586
rect 53170 21534 53182 21586
rect 47070 21522 47122 21534
rect 1934 21474 1986 21486
rect 13246 21474 13298 21486
rect 18510 21474 18562 21486
rect 12674 21422 12686 21474
rect 12738 21422 12750 21474
rect 13794 21422 13806 21474
rect 13858 21422 13870 21474
rect 14690 21422 14702 21474
rect 14754 21422 14766 21474
rect 15586 21422 15598 21474
rect 15650 21422 15662 21474
rect 1934 21410 1986 21422
rect 13246 21410 13298 21422
rect 18510 21410 18562 21422
rect 18734 21474 18786 21486
rect 18734 21410 18786 21422
rect 21422 21474 21474 21486
rect 21422 21410 21474 21422
rect 23774 21474 23826 21486
rect 23774 21410 23826 21422
rect 24222 21474 24274 21486
rect 28030 21474 28082 21486
rect 41246 21474 41298 21486
rect 54462 21474 54514 21486
rect 26562 21422 26574 21474
rect 26626 21422 26638 21474
rect 30034 21422 30046 21474
rect 30098 21422 30110 21474
rect 33842 21422 33854 21474
rect 33906 21422 33918 21474
rect 51650 21422 51662 21474
rect 51714 21422 51726 21474
rect 53330 21422 53342 21474
rect 53394 21422 53406 21474
rect 24222 21410 24274 21422
rect 28030 21410 28082 21422
rect 41246 21410 41298 21422
rect 54462 21410 54514 21422
rect 38446 21362 38498 21374
rect 31266 21310 31278 21362
rect 31330 21310 31342 21362
rect 38446 21298 38498 21310
rect 41582 21362 41634 21374
rect 41582 21298 41634 21310
rect 44718 21362 44770 21374
rect 44718 21298 44770 21310
rect 46734 21362 46786 21374
rect 46734 21298 46786 21310
rect 54350 21362 54402 21374
rect 54350 21298 54402 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 30270 21026 30322 21038
rect 30270 20962 30322 20974
rect 37550 21026 37602 21038
rect 37550 20962 37602 20974
rect 47630 21026 47682 21038
rect 49970 20974 49982 21026
rect 50034 20974 50046 21026
rect 47630 20962 47682 20974
rect 11118 20914 11170 20926
rect 22878 20914 22930 20926
rect 12450 20862 12462 20914
rect 12514 20862 12526 20914
rect 11118 20850 11170 20862
rect 22878 20850 22930 20862
rect 23774 20914 23826 20926
rect 23774 20850 23826 20862
rect 27022 20914 27074 20926
rect 27022 20850 27074 20862
rect 31726 20914 31778 20926
rect 31726 20850 31778 20862
rect 36990 20914 37042 20926
rect 36990 20850 37042 20862
rect 38446 20914 38498 20926
rect 38446 20850 38498 20862
rect 39902 20914 39954 20926
rect 39902 20850 39954 20862
rect 47294 20914 47346 20926
rect 47294 20850 47346 20862
rect 49422 20914 49474 20926
rect 51774 20914 51826 20926
rect 50530 20862 50542 20914
rect 50594 20862 50606 20914
rect 49422 20850 49474 20862
rect 51774 20850 51826 20862
rect 57934 20914 57986 20926
rect 57934 20850 57986 20862
rect 7422 20802 7474 20814
rect 12910 20802 12962 20814
rect 19182 20802 19234 20814
rect 5842 20750 5854 20802
rect 5906 20750 5918 20802
rect 7970 20750 7982 20802
rect 8034 20750 8046 20802
rect 14018 20750 14030 20802
rect 14082 20750 14094 20802
rect 15810 20750 15822 20802
rect 15874 20750 15886 20802
rect 17378 20750 17390 20802
rect 17442 20750 17454 20802
rect 7422 20738 7474 20750
rect 12910 20738 12962 20750
rect 19182 20738 19234 20750
rect 20638 20802 20690 20814
rect 25342 20802 25394 20814
rect 24546 20750 24558 20802
rect 24610 20750 24622 20802
rect 20638 20738 20690 20750
rect 25342 20738 25394 20750
rect 27918 20802 27970 20814
rect 37214 20802 37266 20814
rect 31154 20750 31166 20802
rect 31218 20750 31230 20802
rect 31378 20750 31390 20802
rect 31442 20750 31454 20802
rect 33618 20750 33630 20802
rect 33682 20750 33694 20802
rect 35858 20750 35870 20802
rect 35922 20750 35934 20802
rect 27918 20738 27970 20750
rect 37214 20738 37266 20750
rect 37998 20802 38050 20814
rect 46398 20802 46450 20814
rect 49646 20802 49698 20814
rect 41570 20750 41582 20802
rect 41634 20750 41646 20802
rect 42466 20750 42478 20802
rect 42530 20750 42542 20802
rect 46610 20750 46622 20802
rect 46674 20750 46686 20802
rect 37998 20738 38050 20750
rect 46398 20738 46450 20750
rect 49646 20738 49698 20750
rect 50990 20802 51042 20814
rect 51202 20750 51214 20802
rect 51266 20750 51278 20802
rect 54002 20750 54014 20802
rect 54066 20750 54078 20802
rect 54226 20750 54238 20802
rect 54290 20750 54302 20802
rect 55570 20750 55582 20802
rect 55634 20750 55646 20802
rect 50990 20738 51042 20750
rect 11566 20690 11618 20702
rect 20750 20690 20802 20702
rect 14466 20638 14478 20690
rect 14530 20638 14542 20690
rect 15922 20638 15934 20690
rect 15986 20638 15998 20690
rect 17154 20638 17166 20690
rect 17218 20638 17230 20690
rect 19730 20638 19742 20690
rect 19794 20638 19806 20690
rect 20402 20638 20414 20690
rect 20466 20638 20478 20690
rect 11566 20626 11618 20638
rect 20750 20626 20802 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 21534 20690 21586 20702
rect 21534 20626 21586 20638
rect 21870 20690 21922 20702
rect 21870 20626 21922 20638
rect 22430 20690 22482 20702
rect 25454 20690 25506 20702
rect 24770 20638 24782 20690
rect 24834 20638 24846 20690
rect 22430 20626 22482 20638
rect 25454 20626 25506 20638
rect 25678 20690 25730 20702
rect 25678 20626 25730 20638
rect 30158 20690 30210 20702
rect 30158 20626 30210 20638
rect 31614 20690 31666 20702
rect 36094 20690 36146 20702
rect 33282 20638 33294 20690
rect 33346 20638 33358 20690
rect 35074 20638 35086 20690
rect 35138 20638 35150 20690
rect 31614 20626 31666 20638
rect 36094 20626 36146 20638
rect 40014 20690 40066 20702
rect 40014 20626 40066 20638
rect 40238 20690 40290 20702
rect 40238 20626 40290 20638
rect 40462 20690 40514 20702
rect 40462 20626 40514 20638
rect 40574 20690 40626 20702
rect 45390 20690 45442 20702
rect 41682 20638 41694 20690
rect 41746 20638 41758 20690
rect 40574 20626 40626 20638
rect 45390 20626 45442 20638
rect 47742 20690 47794 20702
rect 47742 20626 47794 20638
rect 50318 20690 50370 20702
rect 50318 20626 50370 20638
rect 54462 20690 54514 20702
rect 54462 20626 54514 20638
rect 54798 20690 54850 20702
rect 54798 20626 54850 20638
rect 55134 20690 55186 20702
rect 55134 20626 55186 20638
rect 6078 20578 6130 20590
rect 6078 20514 6130 20526
rect 6414 20578 6466 20590
rect 10670 20578 10722 20590
rect 6738 20526 6750 20578
rect 6802 20526 6814 20578
rect 7074 20526 7086 20578
rect 7138 20526 7150 20578
rect 7746 20526 7758 20578
rect 7810 20526 7822 20578
rect 6414 20514 6466 20526
rect 10670 20514 10722 20526
rect 12014 20578 12066 20590
rect 12014 20514 12066 20526
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 18622 20578 18674 20590
rect 18622 20514 18674 20526
rect 21758 20578 21810 20590
rect 21758 20514 21810 20526
rect 22094 20578 22146 20590
rect 22094 20514 22146 20526
rect 22318 20578 22370 20590
rect 22318 20514 22370 20526
rect 23326 20578 23378 20590
rect 23326 20514 23378 20526
rect 26126 20578 26178 20590
rect 26126 20514 26178 20526
rect 26574 20578 26626 20590
rect 26574 20514 26626 20526
rect 27358 20578 27410 20590
rect 27358 20514 27410 20526
rect 28366 20578 28418 20590
rect 28366 20514 28418 20526
rect 29374 20578 29426 20590
rect 29374 20514 29426 20526
rect 29934 20578 29986 20590
rect 29934 20514 29986 20526
rect 30270 20578 30322 20590
rect 30270 20514 30322 20526
rect 31838 20578 31890 20590
rect 31838 20514 31890 20526
rect 32846 20578 32898 20590
rect 32846 20514 32898 20526
rect 39790 20578 39842 20590
rect 44830 20578 44882 20590
rect 42466 20526 42478 20578
rect 42530 20526 42542 20578
rect 39790 20514 39842 20526
rect 44830 20514 44882 20526
rect 50542 20578 50594 20590
rect 50542 20514 50594 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 14478 20242 14530 20254
rect 27582 20242 27634 20254
rect 21074 20190 21086 20242
rect 21138 20190 21150 20242
rect 14478 20178 14530 20190
rect 27582 20178 27634 20190
rect 16830 20130 16882 20142
rect 8082 20078 8094 20130
rect 8146 20078 8158 20130
rect 8642 20078 8654 20130
rect 8706 20078 8718 20130
rect 12338 20078 12350 20130
rect 12402 20078 12414 20130
rect 16830 20066 16882 20078
rect 18398 20130 18450 20142
rect 27134 20130 27186 20142
rect 35870 20130 35922 20142
rect 37438 20130 37490 20142
rect 19058 20078 19070 20130
rect 19122 20078 19134 20130
rect 19506 20078 19518 20130
rect 19570 20078 19582 20130
rect 24322 20078 24334 20130
rect 24386 20078 24398 20130
rect 34066 20078 34078 20130
rect 34130 20078 34142 20130
rect 36530 20078 36542 20130
rect 36594 20078 36606 20130
rect 18398 20066 18450 20078
rect 27134 20066 27186 20078
rect 35870 20066 35922 20078
rect 37438 20066 37490 20078
rect 7086 20018 7138 20030
rect 6402 19966 6414 20018
rect 6466 19966 6478 20018
rect 7086 19954 7138 19966
rect 7310 20018 7362 20030
rect 11342 20018 11394 20030
rect 15486 20018 15538 20030
rect 7970 19966 7982 20018
rect 8034 19966 8046 20018
rect 9986 19966 9998 20018
rect 10050 19966 10062 20018
rect 13122 19966 13134 20018
rect 13186 19966 13198 20018
rect 14578 19966 14590 20018
rect 14642 19966 14654 20018
rect 7310 19954 7362 19966
rect 11342 19954 11394 19966
rect 15486 19954 15538 19966
rect 15710 20018 15762 20030
rect 16942 20018 16994 20030
rect 18734 20018 18786 20030
rect 25342 20018 25394 20030
rect 16370 19966 16382 20018
rect 16434 19966 16446 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 17714 19966 17726 20018
rect 17778 19966 17790 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 21186 19966 21198 20018
rect 21250 19966 21262 20018
rect 21522 19966 21534 20018
rect 21586 19966 21598 20018
rect 23314 19966 23326 20018
rect 23378 19966 23390 20018
rect 24098 19966 24110 20018
rect 24162 19966 24174 20018
rect 15710 19954 15762 19966
rect 16942 19954 16994 19966
rect 18734 19954 18786 19966
rect 25342 19954 25394 19966
rect 25678 20018 25730 20030
rect 25678 19954 25730 19966
rect 26238 20018 26290 20030
rect 26238 19954 26290 19966
rect 29038 20018 29090 20030
rect 29038 19954 29090 19966
rect 29262 20018 29314 20030
rect 29262 19954 29314 19966
rect 29710 20018 29762 20030
rect 29710 19954 29762 19966
rect 30382 20018 30434 20030
rect 30382 19954 30434 19966
rect 32398 20018 32450 20030
rect 32398 19954 32450 19966
rect 33518 20018 33570 20030
rect 33518 19954 33570 19966
rect 33742 20018 33794 20030
rect 33742 19954 33794 19966
rect 35198 20018 35250 20030
rect 35198 19954 35250 19966
rect 35646 20018 35698 20030
rect 37998 20018 38050 20030
rect 41582 20018 41634 20030
rect 36306 19966 36318 20018
rect 36370 19966 36382 20018
rect 38210 19966 38222 20018
rect 38274 19966 38286 20018
rect 35646 19954 35698 19966
rect 37998 19954 38050 19966
rect 41582 19954 41634 19966
rect 41918 20018 41970 20030
rect 41918 19954 41970 19966
rect 42142 20018 42194 20030
rect 42142 19954 42194 19966
rect 10558 19906 10610 19918
rect 6066 19854 6078 19906
rect 6130 19854 6142 19906
rect 9650 19854 9662 19906
rect 9714 19854 9726 19906
rect 10434 19854 10446 19906
rect 10498 19854 10510 19906
rect 7634 19742 7646 19794
rect 7698 19742 7710 19794
rect 10449 19791 10495 19854
rect 10558 19842 10610 19854
rect 11006 19906 11058 19918
rect 11006 19842 11058 19854
rect 11902 19906 11954 19918
rect 23774 19906 23826 19918
rect 26798 19906 26850 19918
rect 18050 19854 18062 19906
rect 18114 19854 18126 19906
rect 23986 19854 23998 19906
rect 24050 19854 24062 19906
rect 11902 19842 11954 19854
rect 23774 19842 23826 19854
rect 26798 19842 26850 19854
rect 28142 19906 28194 19918
rect 28142 19842 28194 19854
rect 28478 19906 28530 19918
rect 28478 19842 28530 19854
rect 29150 19906 29202 19918
rect 29150 19842 29202 19854
rect 30046 19906 30098 19918
rect 30046 19842 30098 19854
rect 30942 19906 30994 19918
rect 30942 19842 30994 19854
rect 35422 19906 35474 19918
rect 35422 19842 35474 19854
rect 41806 19906 41858 19918
rect 41806 19842 41858 19854
rect 37102 19794 37154 19806
rect 11106 19791 11118 19794
rect 10449 19745 11118 19791
rect 11106 19742 11118 19745
rect 11170 19742 11182 19794
rect 15138 19742 15150 19794
rect 15202 19742 15214 19794
rect 27346 19742 27358 19794
rect 27410 19791 27422 19794
rect 28466 19791 28478 19794
rect 27410 19745 28478 19791
rect 27410 19742 27422 19745
rect 28466 19742 28478 19745
rect 28530 19742 28542 19794
rect 37102 19730 37154 19742
rect 37886 19794 37938 19806
rect 37886 19730 37938 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 21310 19458 21362 19470
rect 14802 19406 14814 19458
rect 14866 19406 14878 19458
rect 19730 19406 19742 19458
rect 19794 19406 19806 19458
rect 21310 19394 21362 19406
rect 21646 19458 21698 19470
rect 21646 19394 21698 19406
rect 24334 19458 24386 19470
rect 41582 19458 41634 19470
rect 30370 19406 30382 19458
rect 30434 19406 30446 19458
rect 34962 19406 34974 19458
rect 35026 19406 35038 19458
rect 24334 19394 24386 19406
rect 41582 19394 41634 19406
rect 41918 19458 41970 19470
rect 41918 19394 41970 19406
rect 21982 19346 22034 19358
rect 17714 19294 17726 19346
rect 17778 19294 17790 19346
rect 20066 19294 20078 19346
rect 20130 19294 20142 19346
rect 21982 19282 22034 19294
rect 27470 19346 27522 19358
rect 27470 19282 27522 19294
rect 28478 19346 28530 19358
rect 35870 19346 35922 19358
rect 30818 19294 30830 19346
rect 30882 19294 30894 19346
rect 31938 19294 31950 19346
rect 32002 19294 32014 19346
rect 28478 19282 28530 19294
rect 35870 19282 35922 19294
rect 46174 19346 46226 19358
rect 46174 19282 46226 19294
rect 47070 19346 47122 19358
rect 47070 19282 47122 19294
rect 51886 19346 51938 19358
rect 51886 19282 51938 19294
rect 9774 19234 9826 19246
rect 5954 19182 5966 19234
rect 6018 19182 6030 19234
rect 6402 19182 6414 19234
rect 6466 19182 6478 19234
rect 8978 19182 8990 19234
rect 9042 19182 9054 19234
rect 9774 19170 9826 19182
rect 10110 19234 10162 19246
rect 17838 19234 17890 19246
rect 26462 19234 26514 19246
rect 10658 19182 10670 19234
rect 10722 19182 10734 19234
rect 11106 19182 11118 19234
rect 11170 19182 11182 19234
rect 13682 19182 13694 19234
rect 13746 19182 13758 19234
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 18834 19182 18846 19234
rect 18898 19182 18910 19234
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 22418 19182 22430 19234
rect 22482 19182 22494 19234
rect 24882 19182 24894 19234
rect 24946 19182 24958 19234
rect 25778 19182 25790 19234
rect 25842 19182 25854 19234
rect 10110 19170 10162 19182
rect 17838 19170 17890 19182
rect 26462 19170 26514 19182
rect 26686 19234 26738 19246
rect 26686 19170 26738 19182
rect 26798 19234 26850 19246
rect 26798 19170 26850 19182
rect 27694 19234 27746 19246
rect 27694 19170 27746 19182
rect 29262 19234 29314 19246
rect 31502 19234 31554 19246
rect 29474 19182 29486 19234
rect 29538 19182 29550 19234
rect 30482 19182 30494 19234
rect 30546 19182 30558 19234
rect 29262 19170 29314 19182
rect 31502 19170 31554 19182
rect 32734 19234 32786 19246
rect 34302 19234 34354 19246
rect 46958 19234 47010 19246
rect 32946 19182 32958 19234
rect 33010 19182 33022 19234
rect 33842 19182 33854 19234
rect 33906 19182 33918 19234
rect 34402 19182 34414 19234
rect 34466 19182 34478 19234
rect 46610 19182 46622 19234
rect 46674 19182 46686 19234
rect 32734 19170 32786 19182
rect 34302 19170 34354 19182
rect 46958 19170 47010 19182
rect 47630 19234 47682 19246
rect 47630 19170 47682 19182
rect 50766 19234 50818 19246
rect 50766 19170 50818 19182
rect 51326 19234 51378 19246
rect 51326 19170 51378 19182
rect 51550 19234 51602 19246
rect 53218 19182 53230 19234
rect 53282 19182 53294 19234
rect 53554 19182 53566 19234
rect 53618 19182 53630 19234
rect 51550 19170 51602 19182
rect 19294 19122 19346 19134
rect 7410 19070 7422 19122
rect 7474 19070 7486 19122
rect 9202 19070 9214 19122
rect 9266 19070 9278 19122
rect 12114 19070 12126 19122
rect 12178 19070 12190 19122
rect 13570 19070 13582 19122
rect 13634 19070 13646 19122
rect 16034 19070 16046 19122
rect 16098 19070 16110 19122
rect 19294 19058 19346 19070
rect 21534 19122 21586 19134
rect 21534 19058 21586 19070
rect 27134 19122 27186 19134
rect 52882 19070 52894 19122
rect 52946 19070 52958 19122
rect 27134 19058 27186 19070
rect 1710 19010 1762 19022
rect 1710 18946 1762 18958
rect 8654 19010 8706 19022
rect 8654 18946 8706 18958
rect 12910 19010 12962 19022
rect 12910 18946 12962 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 22766 19010 22818 19022
rect 22766 18946 22818 18958
rect 23102 19010 23154 19022
rect 32398 19010 32450 19022
rect 28018 18958 28030 19010
rect 28082 18958 28094 19010
rect 23102 18946 23154 18958
rect 32398 18946 32450 18958
rect 41806 19010 41858 19022
rect 41806 18946 41858 18958
rect 46062 19010 46114 19022
rect 46062 18946 46114 18958
rect 46286 19010 46338 19022
rect 46286 18946 46338 18958
rect 47182 19010 47234 19022
rect 47182 18946 47234 18958
rect 50542 19010 50594 19022
rect 50542 18946 50594 18958
rect 50878 19010 50930 19022
rect 50878 18946 50930 18958
rect 50990 19010 51042 19022
rect 53666 18958 53678 19010
rect 53730 18958 53742 19010
rect 50990 18946 51042 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 7870 18674 7922 18686
rect 7870 18610 7922 18622
rect 8654 18674 8706 18686
rect 8654 18610 8706 18622
rect 11006 18674 11058 18686
rect 11006 18610 11058 18622
rect 18062 18674 18114 18686
rect 18062 18610 18114 18622
rect 18174 18674 18226 18686
rect 18174 18610 18226 18622
rect 24446 18674 24498 18686
rect 24446 18610 24498 18622
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 29598 18674 29650 18686
rect 29598 18610 29650 18622
rect 34526 18674 34578 18686
rect 39554 18622 39566 18674
rect 39618 18622 39630 18674
rect 34526 18610 34578 18622
rect 6750 18562 6802 18574
rect 16942 18562 16994 18574
rect 13122 18510 13134 18562
rect 13186 18510 13198 18562
rect 14466 18510 14478 18562
rect 14530 18510 14542 18562
rect 15250 18510 15262 18562
rect 15314 18510 15326 18562
rect 6750 18498 6802 18510
rect 16942 18498 16994 18510
rect 17838 18562 17890 18574
rect 17838 18498 17890 18510
rect 17950 18562 18002 18574
rect 25678 18562 25730 18574
rect 34414 18562 34466 18574
rect 19170 18510 19182 18562
rect 19234 18510 19246 18562
rect 21186 18510 21198 18562
rect 21250 18510 21262 18562
rect 27682 18510 27694 18562
rect 27746 18510 27758 18562
rect 28354 18510 28366 18562
rect 28418 18510 28430 18562
rect 17950 18498 18002 18510
rect 25678 18498 25730 18510
rect 34414 18498 34466 18510
rect 35198 18562 35250 18574
rect 43374 18562 43426 18574
rect 47070 18562 47122 18574
rect 41234 18510 41246 18562
rect 41298 18510 41310 18562
rect 42578 18510 42590 18562
rect 42642 18510 42654 18562
rect 45714 18510 45726 18562
rect 45778 18510 45790 18562
rect 51986 18510 51998 18562
rect 52050 18510 52062 18562
rect 54226 18510 54238 18562
rect 54290 18510 54302 18562
rect 55122 18510 55134 18562
rect 55186 18510 55198 18562
rect 35198 18498 35250 18510
rect 43374 18498 43426 18510
rect 47070 18498 47122 18510
rect 6974 18450 7026 18462
rect 6974 18386 7026 18398
rect 7198 18450 7250 18462
rect 7198 18386 7250 18398
rect 9102 18450 9154 18462
rect 12798 18450 12850 18462
rect 21758 18450 21810 18462
rect 25454 18450 25506 18462
rect 30270 18450 30322 18462
rect 11778 18398 11790 18450
rect 11842 18398 11854 18450
rect 12338 18398 12350 18450
rect 12402 18398 12414 18450
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 14802 18398 14814 18450
rect 14866 18398 14878 18450
rect 16034 18398 16046 18450
rect 16098 18398 16110 18450
rect 17490 18398 17502 18450
rect 17554 18398 17566 18450
rect 19058 18398 19070 18450
rect 19122 18398 19134 18450
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 23202 18398 23214 18450
rect 23266 18398 23278 18450
rect 26114 18398 26126 18450
rect 26178 18398 26190 18450
rect 27570 18398 27582 18450
rect 27634 18398 27646 18450
rect 28130 18398 28142 18450
rect 28194 18398 28206 18450
rect 29026 18398 29038 18450
rect 29090 18398 29102 18450
rect 9102 18386 9154 18398
rect 12798 18386 12850 18398
rect 21758 18386 21810 18398
rect 25454 18386 25506 18398
rect 30270 18386 30322 18398
rect 30382 18450 30434 18462
rect 33182 18450 33234 18462
rect 34750 18450 34802 18462
rect 30594 18398 30606 18450
rect 30658 18398 30670 18450
rect 33394 18398 33406 18450
rect 33458 18398 33470 18450
rect 30382 18386 30434 18398
rect 33182 18386 33234 18398
rect 34750 18386 34802 18398
rect 35086 18450 35138 18462
rect 35086 18386 35138 18398
rect 35758 18450 35810 18462
rect 38334 18450 38386 18462
rect 37986 18398 37998 18450
rect 38050 18398 38062 18450
rect 35758 18386 35810 18398
rect 38334 18386 38386 18398
rect 38670 18450 38722 18462
rect 42142 18450 42194 18462
rect 39778 18398 39790 18450
rect 39842 18398 39854 18450
rect 41010 18398 41022 18450
rect 41074 18398 41086 18450
rect 38670 18386 38722 18398
rect 42142 18386 42194 18398
rect 42926 18450 42978 18462
rect 42926 18386 42978 18398
rect 43262 18450 43314 18462
rect 43262 18386 43314 18398
rect 43598 18450 43650 18462
rect 43598 18386 43650 18398
rect 43934 18450 43986 18462
rect 44830 18450 44882 18462
rect 47182 18450 47234 18462
rect 44146 18398 44158 18450
rect 44210 18398 44222 18450
rect 45602 18398 45614 18450
rect 45666 18398 45678 18450
rect 46610 18398 46622 18450
rect 46674 18398 46686 18450
rect 43934 18386 43986 18398
rect 44830 18386 44882 18398
rect 47182 18386 47234 18398
rect 47294 18450 47346 18462
rect 47294 18386 47346 18398
rect 47742 18450 47794 18462
rect 49870 18450 49922 18462
rect 48962 18398 48974 18450
rect 49026 18398 49038 18450
rect 51090 18398 51102 18450
rect 51154 18398 51166 18450
rect 52546 18398 52558 18450
rect 52610 18398 52622 18450
rect 53778 18398 53790 18450
rect 53842 18398 53854 18450
rect 55682 18398 55694 18450
rect 55746 18398 55758 18450
rect 47742 18386 47794 18398
rect 49870 18386 49922 18398
rect 9662 18338 9714 18350
rect 9662 18274 9714 18286
rect 10110 18338 10162 18350
rect 18846 18338 18898 18350
rect 10546 18286 10558 18338
rect 10610 18286 10622 18338
rect 11442 18286 11454 18338
rect 11506 18286 11518 18338
rect 13794 18286 13806 18338
rect 13858 18286 13870 18338
rect 10110 18274 10162 18286
rect 18846 18274 18898 18286
rect 23662 18338 23714 18350
rect 23662 18274 23714 18286
rect 26910 18338 26962 18350
rect 26910 18274 26962 18286
rect 31054 18338 31106 18350
rect 31054 18274 31106 18286
rect 31950 18338 32002 18350
rect 31950 18274 32002 18286
rect 39230 18338 39282 18350
rect 51550 18338 51602 18350
rect 45826 18286 45838 18338
rect 45890 18286 45902 18338
rect 49186 18286 49198 18338
rect 49250 18286 49262 18338
rect 50754 18286 50766 18338
rect 50818 18286 50830 18338
rect 39230 18274 39282 18286
rect 51550 18274 51602 18286
rect 7422 18226 7474 18238
rect 7422 18162 7474 18174
rect 14702 18226 14754 18238
rect 14702 18162 14754 18174
rect 24334 18226 24386 18238
rect 32174 18226 32226 18238
rect 35198 18226 35250 18238
rect 29810 18174 29822 18226
rect 29874 18174 29886 18226
rect 32498 18174 32510 18226
rect 32562 18174 32574 18226
rect 33842 18174 33854 18226
rect 33906 18174 33918 18226
rect 24334 18162 24386 18174
rect 32174 18162 32226 18174
rect 35198 18162 35250 18174
rect 41806 18226 41858 18238
rect 41806 18162 41858 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 34302 17890 34354 17902
rect 30482 17838 30494 17890
rect 30546 17838 30558 17890
rect 34302 17826 34354 17838
rect 42814 17890 42866 17902
rect 42814 17826 42866 17838
rect 45502 17890 45554 17902
rect 45502 17826 45554 17838
rect 49198 17890 49250 17902
rect 49198 17826 49250 17838
rect 49534 17890 49586 17902
rect 49534 17826 49586 17838
rect 11902 17778 11954 17790
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 11902 17714 11954 17726
rect 12910 17778 12962 17790
rect 12910 17714 12962 17726
rect 27022 17778 27074 17790
rect 27022 17714 27074 17726
rect 28142 17778 28194 17790
rect 33742 17778 33794 17790
rect 30594 17726 30606 17778
rect 30658 17726 30670 17778
rect 28142 17714 28194 17726
rect 33742 17714 33794 17726
rect 36542 17778 36594 17790
rect 36542 17714 36594 17726
rect 37550 17778 37602 17790
rect 37550 17714 37602 17726
rect 46846 17778 46898 17790
rect 46846 17714 46898 17726
rect 48974 17778 49026 17790
rect 48974 17714 49026 17726
rect 52558 17778 52610 17790
rect 57934 17778 57986 17790
rect 54338 17726 54350 17778
rect 54402 17726 54414 17778
rect 52558 17714 52610 17726
rect 57934 17714 57986 17726
rect 9550 17666 9602 17678
rect 9550 17602 9602 17614
rect 10670 17666 10722 17678
rect 10670 17602 10722 17614
rect 11342 17666 11394 17678
rect 18286 17666 18338 17678
rect 20414 17666 20466 17678
rect 23774 17666 23826 17678
rect 12450 17614 12462 17666
rect 12514 17614 12526 17666
rect 13906 17614 13918 17666
rect 13970 17614 13982 17666
rect 14354 17614 14366 17666
rect 14418 17614 14430 17666
rect 15810 17614 15822 17666
rect 15874 17614 15886 17666
rect 16818 17614 16830 17666
rect 16882 17614 16894 17666
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 21410 17614 21422 17666
rect 21474 17614 21486 17666
rect 11342 17602 11394 17614
rect 18286 17602 18338 17614
rect 20414 17602 20466 17614
rect 23774 17602 23826 17614
rect 24446 17666 24498 17678
rect 24446 17602 24498 17614
rect 25118 17666 25170 17678
rect 33182 17666 33234 17678
rect 29586 17614 29598 17666
rect 29650 17614 29662 17666
rect 30706 17614 30718 17666
rect 30770 17614 30782 17666
rect 25118 17602 25170 17614
rect 33182 17602 33234 17614
rect 35086 17666 35138 17678
rect 38782 17666 38834 17678
rect 37202 17614 37214 17666
rect 37266 17614 37278 17666
rect 35086 17602 35138 17614
rect 38782 17602 38834 17614
rect 39342 17666 39394 17678
rect 41694 17666 41746 17678
rect 50990 17666 51042 17678
rect 40898 17614 40910 17666
rect 40962 17614 40974 17666
rect 45490 17614 45502 17666
rect 45554 17614 45566 17666
rect 46386 17614 46398 17666
rect 46450 17614 46462 17666
rect 50418 17614 50430 17666
rect 50482 17614 50494 17666
rect 39342 17602 39394 17614
rect 41694 17602 41746 17614
rect 50990 17602 51042 17614
rect 52670 17666 52722 17678
rect 54562 17614 54574 17666
rect 54626 17614 54638 17666
rect 55570 17614 55582 17666
rect 55634 17614 55646 17666
rect 52670 17602 52722 17614
rect 18174 17554 18226 17566
rect 22542 17554 22594 17566
rect 17154 17502 17166 17554
rect 17218 17502 17230 17554
rect 21634 17502 21646 17554
rect 21698 17502 21710 17554
rect 21970 17502 21982 17554
rect 22034 17502 22046 17554
rect 18174 17490 18226 17502
rect 22542 17490 22594 17502
rect 23438 17554 23490 17566
rect 31950 17554 32002 17566
rect 24098 17502 24110 17554
rect 24162 17502 24174 17554
rect 23438 17490 23490 17502
rect 31950 17490 32002 17502
rect 34190 17554 34242 17566
rect 34190 17490 34242 17502
rect 34750 17554 34802 17566
rect 34750 17490 34802 17502
rect 34862 17554 34914 17566
rect 34862 17490 34914 17502
rect 37774 17554 37826 17566
rect 38446 17554 38498 17566
rect 37874 17502 37886 17554
rect 37938 17551 37950 17554
rect 38210 17551 38222 17554
rect 37938 17505 38222 17551
rect 37938 17502 37950 17505
rect 38210 17502 38222 17505
rect 38274 17502 38286 17554
rect 37774 17490 37826 17502
rect 38446 17490 38498 17502
rect 39006 17554 39058 17566
rect 42590 17554 42642 17566
rect 41122 17502 41134 17554
rect 41186 17502 41198 17554
rect 39006 17490 39058 17502
rect 42590 17490 42642 17502
rect 42702 17554 42754 17566
rect 42702 17490 42754 17502
rect 45166 17554 45218 17566
rect 45166 17490 45218 17502
rect 51102 17554 51154 17566
rect 55134 17554 55186 17566
rect 52882 17502 52894 17554
rect 52946 17502 52958 17554
rect 53442 17502 53454 17554
rect 53506 17502 53518 17554
rect 51102 17490 51154 17502
rect 55134 17490 55186 17502
rect 1710 17442 1762 17454
rect 1710 17378 1762 17390
rect 7982 17442 8034 17454
rect 7982 17378 8034 17390
rect 8430 17442 8482 17454
rect 8430 17378 8482 17390
rect 8878 17442 8930 17454
rect 8878 17378 8930 17390
rect 9326 17442 9378 17454
rect 9326 17378 9378 17390
rect 11118 17442 11170 17454
rect 11118 17378 11170 17390
rect 13582 17442 13634 17454
rect 13582 17378 13634 17390
rect 16270 17442 16322 17454
rect 22990 17442 23042 17454
rect 25230 17442 25282 17454
rect 20738 17390 20750 17442
rect 20802 17390 20814 17442
rect 24770 17390 24782 17442
rect 24834 17390 24846 17442
rect 16270 17378 16322 17390
rect 22990 17378 23042 17390
rect 25230 17378 25282 17390
rect 25454 17442 25506 17454
rect 25454 17378 25506 17390
rect 26126 17442 26178 17454
rect 26126 17378 26178 17390
rect 26574 17442 26626 17454
rect 26574 17378 26626 17390
rect 27582 17442 27634 17454
rect 27582 17378 27634 17390
rect 28702 17442 28754 17454
rect 28702 17378 28754 17390
rect 29374 17442 29426 17454
rect 29374 17378 29426 17390
rect 31502 17442 31554 17454
rect 31502 17378 31554 17390
rect 32510 17442 32562 17454
rect 32510 17378 32562 17390
rect 32958 17442 33010 17454
rect 32958 17378 33010 17390
rect 33630 17442 33682 17454
rect 33630 17378 33682 17390
rect 33854 17442 33906 17454
rect 33854 17378 33906 17390
rect 34302 17442 34354 17454
rect 34302 17378 34354 17390
rect 35982 17442 36034 17454
rect 35982 17378 36034 17390
rect 38894 17442 38946 17454
rect 40126 17442 40178 17454
rect 39666 17390 39678 17442
rect 39730 17390 39742 17442
rect 38894 17378 38946 17390
rect 40126 17378 40178 17390
rect 42030 17442 42082 17454
rect 42030 17378 42082 17390
rect 46734 17442 46786 17454
rect 46734 17378 46786 17390
rect 46958 17442 47010 17454
rect 47630 17442 47682 17454
rect 47282 17390 47294 17442
rect 47346 17390 47358 17442
rect 46958 17378 47010 17390
rect 47630 17378 47682 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 5406 17106 5458 17118
rect 5406 17042 5458 17054
rect 7310 17106 7362 17118
rect 7310 17042 7362 17054
rect 9886 17106 9938 17118
rect 9886 17042 9938 17054
rect 17838 17106 17890 17118
rect 17838 17042 17890 17054
rect 26910 17106 26962 17118
rect 26910 17042 26962 17054
rect 27918 17106 27970 17118
rect 27918 17042 27970 17054
rect 28142 17106 28194 17118
rect 28142 17042 28194 17054
rect 32622 17106 32674 17118
rect 32622 17042 32674 17054
rect 33070 17106 33122 17118
rect 39678 17106 39730 17118
rect 33394 17054 33406 17106
rect 33458 17054 33470 17106
rect 33070 17042 33122 17054
rect 39678 17042 39730 17054
rect 39902 17106 39954 17118
rect 53230 17106 53282 17118
rect 47058 17054 47070 17106
rect 47122 17054 47134 17106
rect 39902 17042 39954 17054
rect 53230 17042 53282 17054
rect 54350 17106 54402 17118
rect 54350 17042 54402 17054
rect 54462 17106 54514 17118
rect 54462 17042 54514 17054
rect 55246 17106 55298 17118
rect 55246 17042 55298 17054
rect 7646 16994 7698 17006
rect 6066 16942 6078 16994
rect 6130 16942 6142 16994
rect 6514 16942 6526 16994
rect 6578 16942 6590 16994
rect 7646 16930 7698 16942
rect 8990 16994 9042 17006
rect 23774 16994 23826 17006
rect 34190 16994 34242 17006
rect 10770 16942 10782 16994
rect 10834 16942 10846 16994
rect 12002 16942 12014 16994
rect 12066 16942 12078 16994
rect 25890 16942 25902 16994
rect 25954 16942 25966 16994
rect 8990 16930 9042 16942
rect 23774 16930 23826 16942
rect 34190 16930 34242 16942
rect 34414 16994 34466 17006
rect 34414 16930 34466 16942
rect 34526 16994 34578 17006
rect 34526 16930 34578 16942
rect 34974 16994 35026 17006
rect 34974 16930 35026 16942
rect 35086 16994 35138 17006
rect 46286 16994 46338 17006
rect 38210 16942 38222 16994
rect 38274 16942 38286 16994
rect 41458 16942 41470 16994
rect 41522 16942 41534 16994
rect 45042 16942 45054 16994
rect 45106 16942 45118 16994
rect 35086 16930 35138 16942
rect 46286 16930 46338 16942
rect 6974 16882 7026 16894
rect 6974 16818 7026 16830
rect 8430 16882 8482 16894
rect 13358 16882 13410 16894
rect 18174 16882 18226 16894
rect 19854 16882 19906 16894
rect 27470 16882 27522 16894
rect 11554 16830 11566 16882
rect 11618 16830 11630 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 18946 16830 18958 16882
rect 19010 16830 19022 16882
rect 20290 16830 20302 16882
rect 20354 16830 20366 16882
rect 23202 16830 23214 16882
rect 23266 16830 23278 16882
rect 24322 16830 24334 16882
rect 24386 16830 24398 16882
rect 25554 16830 25566 16882
rect 25618 16830 25630 16882
rect 26338 16830 26350 16882
rect 26402 16830 26414 16882
rect 8430 16818 8482 16830
rect 13358 16818 13410 16830
rect 18174 16818 18226 16830
rect 19854 16818 19906 16830
rect 27470 16818 27522 16830
rect 27806 16882 27858 16894
rect 29150 16882 29202 16894
rect 35310 16882 35362 16894
rect 28354 16830 28366 16882
rect 28418 16830 28430 16882
rect 31378 16830 31390 16882
rect 31442 16830 31454 16882
rect 33954 16830 33966 16882
rect 34018 16830 34030 16882
rect 27806 16818 27858 16830
rect 29150 16818 29202 16830
rect 35310 16818 35362 16830
rect 37550 16882 37602 16894
rect 39566 16882 39618 16894
rect 46734 16882 46786 16894
rect 38322 16830 38334 16882
rect 38386 16830 38398 16882
rect 39106 16830 39118 16882
rect 39170 16830 39182 16882
rect 41346 16830 41358 16882
rect 41410 16830 41422 16882
rect 44594 16830 44606 16882
rect 44658 16830 44670 16882
rect 45490 16830 45502 16882
rect 45554 16830 45566 16882
rect 37550 16818 37602 16830
rect 39566 16818 39618 16830
rect 46734 16818 46786 16830
rect 53566 16882 53618 16894
rect 55010 16830 55022 16882
rect 55074 16830 55086 16882
rect 53566 16818 53618 16830
rect 5742 16770 5794 16782
rect 23886 16770 23938 16782
rect 36990 16770 37042 16782
rect 46062 16770 46114 16782
rect 13794 16718 13806 16770
rect 13858 16718 13870 16770
rect 16146 16718 16158 16770
rect 16210 16718 16222 16770
rect 22418 16718 22430 16770
rect 22482 16718 22494 16770
rect 25666 16718 25678 16770
rect 25730 16718 25742 16770
rect 29474 16718 29486 16770
rect 29538 16718 29550 16770
rect 31826 16718 31838 16770
rect 31890 16718 31902 16770
rect 38770 16718 38782 16770
rect 38834 16718 38846 16770
rect 41794 16718 41806 16770
rect 41858 16718 41870 16770
rect 45266 16718 45278 16770
rect 45330 16718 45342 16770
rect 46386 16718 46398 16770
rect 46450 16718 46462 16770
rect 53330 16718 53342 16770
rect 53394 16718 53406 16770
rect 5742 16706 5794 16718
rect 23886 16706 23938 16718
rect 36990 16706 37042 16718
rect 46062 16706 46114 16718
rect 7758 16658 7810 16670
rect 7758 16594 7810 16606
rect 10334 16658 10386 16670
rect 24110 16658 24162 16670
rect 22754 16606 22766 16658
rect 22818 16606 22830 16658
rect 10334 16594 10386 16606
rect 24110 16594 24162 16606
rect 54238 16658 54290 16670
rect 54238 16594 54290 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 7870 16322 7922 16334
rect 7870 16258 7922 16270
rect 8206 16322 8258 16334
rect 8206 16258 8258 16270
rect 9998 16322 10050 16334
rect 9998 16258 10050 16270
rect 10222 16322 10274 16334
rect 31390 16322 31442 16334
rect 20066 16270 20078 16322
rect 20130 16270 20142 16322
rect 10222 16258 10274 16270
rect 31390 16258 31442 16270
rect 37774 16322 37826 16334
rect 37774 16258 37826 16270
rect 42366 16322 42418 16334
rect 42366 16258 42418 16270
rect 45166 16322 45218 16334
rect 52098 16270 52110 16322
rect 52162 16270 52174 16322
rect 45166 16258 45218 16270
rect 5854 16210 5906 16222
rect 5854 16146 5906 16158
rect 11566 16210 11618 16222
rect 11566 16146 11618 16158
rect 12014 16210 12066 16222
rect 12014 16146 12066 16158
rect 12574 16210 12626 16222
rect 12574 16146 12626 16158
rect 12910 16210 12962 16222
rect 21646 16210 21698 16222
rect 32958 16210 33010 16222
rect 14130 16158 14142 16210
rect 14194 16158 14206 16210
rect 26562 16158 26574 16210
rect 26626 16158 26638 16210
rect 27906 16158 27918 16210
rect 27970 16158 27982 16210
rect 12910 16146 12962 16158
rect 21646 16146 21698 16158
rect 32958 16146 33010 16158
rect 34302 16210 34354 16222
rect 34302 16146 34354 16158
rect 42142 16210 42194 16222
rect 49534 16210 49586 16222
rect 47170 16158 47182 16210
rect 47234 16158 47246 16210
rect 42142 16146 42194 16158
rect 49534 16146 49586 16158
rect 51774 16210 51826 16222
rect 53678 16210 53730 16222
rect 52994 16158 53006 16210
rect 53058 16158 53070 16210
rect 51774 16146 51826 16158
rect 53678 16146 53730 16158
rect 6414 16098 6466 16110
rect 6414 16034 6466 16046
rect 7086 16098 7138 16110
rect 7086 16034 7138 16046
rect 8542 16098 8594 16110
rect 8542 16034 8594 16046
rect 9102 16098 9154 16110
rect 9102 16034 9154 16046
rect 9886 16098 9938 16110
rect 33406 16098 33458 16110
rect 47518 16098 47570 16110
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 14578 16046 14590 16098
rect 14642 16046 14654 16098
rect 15362 16046 15374 16098
rect 15426 16046 15438 16098
rect 15810 16046 15822 16098
rect 15874 16046 15886 16098
rect 18162 16046 18174 16098
rect 18226 16046 18238 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 19954 16046 19966 16098
rect 20018 16046 20030 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 21746 16046 21758 16098
rect 21810 16046 21822 16098
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 24546 16046 24558 16098
rect 24610 16046 24622 16098
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 26226 16046 26238 16098
rect 26290 16046 26302 16098
rect 26898 16046 26910 16098
rect 26962 16046 26974 16098
rect 27458 16046 27470 16098
rect 27522 16046 27534 16098
rect 29810 16046 29822 16098
rect 29874 16046 29886 16098
rect 30818 16046 30830 16098
rect 30882 16046 30894 16098
rect 33730 16046 33742 16098
rect 33794 16046 33806 16098
rect 37762 16046 37774 16098
rect 37826 16046 37838 16098
rect 39554 16046 39566 16098
rect 39618 16046 39630 16098
rect 39890 16046 39902 16098
rect 39954 16046 39966 16098
rect 41458 16046 41470 16098
rect 41522 16046 41534 16098
rect 43922 16046 43934 16098
rect 43986 16046 43998 16098
rect 45154 16046 45166 16098
rect 45218 16046 45230 16098
rect 46162 16046 46174 16098
rect 46226 16046 46238 16098
rect 46946 16046 46958 16098
rect 47010 16046 47022 16098
rect 9886 16034 9938 16046
rect 33406 16034 33458 16046
rect 47518 16034 47570 16046
rect 47966 16098 48018 16110
rect 47966 16034 48018 16046
rect 48190 16098 48242 16110
rect 48190 16034 48242 16046
rect 51550 16098 51602 16110
rect 52882 16046 52894 16098
rect 52946 16046 52958 16098
rect 51550 16034 51602 16046
rect 6974 15986 7026 15998
rect 6974 15922 7026 15934
rect 7646 15986 7698 15998
rect 22094 15986 22146 15998
rect 37438 15986 37490 15998
rect 44830 15986 44882 15998
rect 14914 15934 14926 15986
rect 14978 15934 14990 15986
rect 18386 15934 18398 15986
rect 18450 15934 18462 15986
rect 27570 15934 27582 15986
rect 27634 15934 27646 15986
rect 30034 15934 30046 15986
rect 30098 15934 30110 15986
rect 30930 15934 30942 15986
rect 30994 15934 31006 15986
rect 38546 15934 38558 15986
rect 38610 15934 38622 15986
rect 44146 15934 44158 15986
rect 44210 15934 44222 15986
rect 47058 15934 47070 15986
rect 47122 15934 47134 15986
rect 7646 15922 7698 15934
rect 22094 15922 22146 15934
rect 37438 15922 37490 15934
rect 44830 15922 44882 15934
rect 6750 15874 6802 15886
rect 6066 15822 6078 15874
rect 6130 15822 6142 15874
rect 6750 15810 6802 15822
rect 10670 15874 10722 15886
rect 10670 15810 10722 15822
rect 18846 15874 18898 15886
rect 18846 15810 18898 15822
rect 21310 15874 21362 15886
rect 21310 15810 21362 15822
rect 21534 15874 21586 15886
rect 21534 15810 21586 15822
rect 28590 15874 28642 15886
rect 28590 15810 28642 15822
rect 36542 15874 36594 15886
rect 36542 15810 36594 15822
rect 37102 15874 37154 15886
rect 48078 15874 48130 15886
rect 39330 15822 39342 15874
rect 39394 15822 39406 15874
rect 42690 15822 42702 15874
rect 42754 15822 42766 15874
rect 37102 15810 37154 15822
rect 48078 15810 48130 15822
rect 49646 15874 49698 15886
rect 49646 15810 49698 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 10782 15538 10834 15550
rect 10782 15474 10834 15486
rect 15822 15538 15874 15550
rect 25342 15538 25394 15550
rect 28814 15538 28866 15550
rect 23426 15486 23438 15538
rect 23490 15486 23502 15538
rect 26338 15486 26350 15538
rect 26402 15486 26414 15538
rect 15822 15474 15874 15486
rect 25342 15474 25394 15486
rect 28814 15474 28866 15486
rect 33630 15538 33682 15550
rect 33630 15474 33682 15486
rect 34638 15538 34690 15550
rect 34638 15474 34690 15486
rect 35870 15538 35922 15550
rect 37886 15538 37938 15550
rect 37090 15486 37102 15538
rect 37154 15486 37166 15538
rect 35870 15474 35922 15486
rect 37886 15474 37938 15486
rect 39790 15538 39842 15550
rect 39790 15474 39842 15486
rect 51102 15538 51154 15550
rect 51102 15474 51154 15486
rect 51214 15538 51266 15550
rect 51214 15474 51266 15486
rect 52782 15538 52834 15550
rect 52782 15474 52834 15486
rect 9550 15426 9602 15438
rect 9550 15362 9602 15374
rect 10110 15426 10162 15438
rect 16830 15426 16882 15438
rect 10434 15374 10446 15426
rect 10498 15374 10510 15426
rect 11778 15374 11790 15426
rect 11842 15374 11854 15426
rect 12674 15374 12686 15426
rect 12738 15374 12750 15426
rect 16258 15374 16270 15426
rect 16322 15374 16334 15426
rect 10110 15362 10162 15374
rect 16830 15362 16882 15374
rect 19854 15426 19906 15438
rect 28254 15426 28306 15438
rect 20402 15374 20414 15426
rect 20466 15374 20478 15426
rect 21746 15374 21758 15426
rect 21810 15374 21822 15426
rect 22530 15374 22542 15426
rect 22594 15374 22606 15426
rect 25778 15374 25790 15426
rect 25842 15374 25854 15426
rect 27346 15374 27358 15426
rect 27410 15374 27422 15426
rect 19854 15362 19906 15374
rect 28254 15362 28306 15374
rect 29150 15426 29202 15438
rect 29150 15362 29202 15374
rect 30046 15426 30098 15438
rect 30046 15362 30098 15374
rect 30158 15426 30210 15438
rect 30158 15362 30210 15374
rect 31614 15426 31666 15438
rect 31614 15362 31666 15374
rect 32062 15426 32114 15438
rect 32062 15362 32114 15374
rect 33742 15426 33794 15438
rect 33742 15362 33794 15374
rect 34302 15426 34354 15438
rect 34302 15362 34354 15374
rect 34414 15426 34466 15438
rect 42030 15426 42082 15438
rect 36418 15374 36430 15426
rect 36482 15374 36494 15426
rect 38322 15374 38334 15426
rect 38386 15374 38398 15426
rect 34414 15362 34466 15374
rect 42030 15362 42082 15374
rect 43374 15426 43426 15438
rect 43374 15362 43426 15374
rect 52670 15426 52722 15438
rect 52670 15362 52722 15374
rect 5630 15314 5682 15326
rect 15262 15314 15314 15326
rect 6514 15262 6526 15314
rect 6578 15262 6590 15314
rect 8754 15262 8766 15314
rect 8818 15262 8830 15314
rect 12450 15262 12462 15314
rect 12514 15262 12526 15314
rect 12786 15262 12798 15314
rect 12850 15262 12862 15314
rect 5630 15250 5682 15262
rect 15262 15250 15314 15262
rect 16606 15314 16658 15326
rect 17950 15314 18002 15326
rect 19630 15314 19682 15326
rect 17602 15262 17614 15314
rect 17666 15262 17678 15314
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 16606 15250 16658 15262
rect 17950 15250 18002 15262
rect 19630 15250 19682 15262
rect 19966 15314 20018 15326
rect 26798 15314 26850 15326
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 22754 15262 22766 15314
rect 22818 15262 22830 15314
rect 24322 15262 24334 15314
rect 24386 15262 24398 15314
rect 25666 15262 25678 15314
rect 25730 15262 25742 15314
rect 19966 15250 20018 15262
rect 26798 15250 26850 15262
rect 27694 15314 27746 15326
rect 31166 15314 31218 15326
rect 33182 15314 33234 15326
rect 29362 15262 29374 15314
rect 29426 15262 29438 15314
rect 30370 15262 30382 15314
rect 30434 15262 30446 15314
rect 31826 15262 31838 15314
rect 31890 15262 31902 15314
rect 27694 15250 27746 15262
rect 31166 15250 31218 15262
rect 33182 15250 33234 15262
rect 33854 15314 33906 15326
rect 33854 15250 33906 15262
rect 34974 15314 35026 15326
rect 49086 15314 49138 15326
rect 50542 15314 50594 15326
rect 36082 15262 36094 15314
rect 36146 15262 36158 15314
rect 36978 15262 36990 15314
rect 37042 15262 37054 15314
rect 38210 15262 38222 15314
rect 38274 15262 38286 15314
rect 39218 15262 39230 15314
rect 39282 15262 39294 15314
rect 42466 15262 42478 15314
rect 42530 15262 42542 15314
rect 49410 15262 49422 15314
rect 49474 15262 49486 15314
rect 34974 15250 35026 15262
rect 49086 15250 49138 15262
rect 50542 15250 50594 15262
rect 50990 15314 51042 15326
rect 53554 15262 53566 15314
rect 53618 15262 53630 15314
rect 50990 15250 51042 15262
rect 6078 15202 6130 15214
rect 15038 15202 15090 15214
rect 24558 15202 24610 15214
rect 6626 15150 6638 15202
rect 6690 15150 6702 15202
rect 14466 15150 14478 15202
rect 14530 15150 14542 15202
rect 18610 15150 18622 15202
rect 18674 15150 18686 15202
rect 21746 15150 21758 15202
rect 21810 15150 21822 15202
rect 6078 15138 6130 15150
rect 15038 15138 15090 15150
rect 24558 15138 24610 15150
rect 24670 15202 24722 15214
rect 40238 15202 40290 15214
rect 32162 15150 32174 15202
rect 32226 15150 32238 15202
rect 38658 15150 38670 15202
rect 38722 15150 38734 15202
rect 24670 15138 24722 15150
rect 40238 15138 40290 15150
rect 41246 15202 41298 15214
rect 45950 15202 46002 15214
rect 42914 15150 42926 15202
rect 42978 15150 42990 15202
rect 41246 15138 41298 15150
rect 45950 15138 46002 15150
rect 48862 15202 48914 15214
rect 48862 15138 48914 15150
rect 49758 15202 49810 15214
rect 49758 15138 49810 15150
rect 49982 15202 50034 15214
rect 49982 15138 50034 15150
rect 52894 15202 52946 15214
rect 54238 15202 54290 15214
rect 53330 15150 53342 15202
rect 53394 15150 53406 15202
rect 52894 15138 52946 15150
rect 54238 15138 54290 15150
rect 31278 15090 31330 15102
rect 8306 15038 8318 15090
rect 8370 15038 8382 15090
rect 14690 15038 14702 15090
rect 14754 15038 14766 15090
rect 18722 15038 18734 15090
rect 18786 15038 18798 15090
rect 31278 15026 31330 15038
rect 50318 15090 50370 15102
rect 50318 15026 50370 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 7646 14754 7698 14766
rect 7646 14690 7698 14702
rect 25790 14754 25842 14766
rect 37998 14754 38050 14766
rect 33282 14702 33294 14754
rect 33346 14702 33358 14754
rect 25790 14690 25842 14702
rect 37998 14690 38050 14702
rect 57934 14754 57986 14766
rect 57934 14690 57986 14702
rect 11342 14642 11394 14654
rect 7298 14590 7310 14642
rect 7362 14639 7374 14642
rect 7522 14639 7534 14642
rect 7362 14593 7534 14639
rect 7362 14590 7374 14593
rect 7522 14590 7534 14593
rect 7586 14590 7598 14642
rect 8306 14590 8318 14642
rect 8370 14590 8382 14642
rect 11342 14578 11394 14590
rect 11790 14642 11842 14654
rect 15374 14642 15426 14654
rect 28590 14642 28642 14654
rect 12786 14590 12798 14642
rect 12850 14590 12862 14642
rect 14578 14590 14590 14642
rect 14642 14590 14654 14642
rect 16706 14590 16718 14642
rect 16770 14590 16782 14642
rect 23762 14590 23774 14642
rect 23826 14590 23838 14642
rect 26114 14590 26126 14642
rect 26178 14590 26190 14642
rect 11790 14578 11842 14590
rect 15374 14578 15426 14590
rect 28590 14578 28642 14590
rect 33854 14642 33906 14654
rect 33854 14578 33906 14590
rect 43598 14642 43650 14654
rect 46398 14642 46450 14654
rect 45490 14590 45502 14642
rect 45554 14590 45566 14642
rect 49074 14590 49086 14642
rect 49138 14590 49150 14642
rect 43598 14578 43650 14590
rect 46398 14578 46450 14590
rect 6190 14530 6242 14542
rect 6190 14466 6242 14478
rect 6638 14530 6690 14542
rect 9214 14530 9266 14542
rect 21198 14530 21250 14542
rect 7746 14478 7758 14530
rect 7810 14478 7822 14530
rect 8530 14478 8542 14530
rect 8594 14478 8606 14530
rect 9538 14478 9550 14530
rect 9602 14478 9614 14530
rect 10210 14478 10222 14530
rect 10274 14478 10286 14530
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 13010 14478 13022 14530
rect 13074 14478 13086 14530
rect 13458 14478 13470 14530
rect 13522 14478 13534 14530
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 18834 14478 18846 14530
rect 18898 14478 18910 14530
rect 19394 14478 19406 14530
rect 19458 14478 19470 14530
rect 19730 14478 19742 14530
rect 19794 14478 19806 14530
rect 6638 14466 6690 14478
rect 9214 14466 9266 14478
rect 21198 14466 21250 14478
rect 21534 14530 21586 14542
rect 27470 14530 27522 14542
rect 22306 14478 22318 14530
rect 22370 14478 22382 14530
rect 22978 14478 22990 14530
rect 23042 14478 23054 14530
rect 23986 14478 23998 14530
rect 24050 14478 24062 14530
rect 24434 14478 24446 14530
rect 24498 14478 24510 14530
rect 21534 14466 21586 14478
rect 27470 14466 27522 14478
rect 29710 14530 29762 14542
rect 31950 14530 32002 14542
rect 33630 14530 33682 14542
rect 30146 14478 30158 14530
rect 30210 14478 30222 14530
rect 31266 14478 31278 14530
rect 31330 14478 31342 14530
rect 32610 14478 32622 14530
rect 32674 14478 32686 14530
rect 29710 14466 29762 14478
rect 31950 14466 32002 14478
rect 33630 14466 33682 14478
rect 33966 14530 34018 14542
rect 33966 14466 34018 14478
rect 34190 14530 34242 14542
rect 34190 14466 34242 14478
rect 36430 14530 36482 14542
rect 41022 14530 41074 14542
rect 46286 14530 46338 14542
rect 38658 14478 38670 14530
rect 38722 14478 38734 14530
rect 40226 14478 40238 14530
rect 40290 14478 40302 14530
rect 41906 14478 41918 14530
rect 41970 14478 41982 14530
rect 45378 14478 45390 14530
rect 45442 14478 45454 14530
rect 36430 14466 36482 14478
rect 41022 14466 41074 14478
rect 46286 14466 46338 14478
rect 47182 14530 47234 14542
rect 54238 14530 54290 14542
rect 47394 14478 47406 14530
rect 47458 14478 47470 14530
rect 48738 14478 48750 14530
rect 48802 14478 48814 14530
rect 50082 14478 50094 14530
rect 50146 14478 50158 14530
rect 55570 14478 55582 14530
rect 55634 14478 55646 14530
rect 47182 14466 47234 14478
rect 54238 14466 54290 14478
rect 6414 14418 6466 14430
rect 6414 14354 6466 14366
rect 9774 14418 9826 14430
rect 21422 14418 21474 14430
rect 24894 14418 24946 14430
rect 10434 14366 10446 14418
rect 10498 14366 10510 14418
rect 10658 14366 10670 14418
rect 10722 14366 10734 14418
rect 16258 14366 16270 14418
rect 16322 14366 16334 14418
rect 19842 14366 19854 14418
rect 19906 14366 19918 14418
rect 21858 14366 21870 14418
rect 21922 14366 21934 14418
rect 23650 14366 23662 14418
rect 23714 14366 23726 14418
rect 9774 14354 9826 14366
rect 21422 14354 21474 14366
rect 24894 14354 24946 14366
rect 25454 14418 25506 14430
rect 27694 14418 27746 14430
rect 26562 14366 26574 14418
rect 26626 14366 26638 14418
rect 27122 14366 27134 14418
rect 27186 14366 27198 14418
rect 25454 14354 25506 14366
rect 27694 14354 27746 14366
rect 27918 14418 27970 14430
rect 36094 14418 36146 14430
rect 34626 14366 34638 14418
rect 34690 14366 34702 14418
rect 27918 14354 27970 14366
rect 36094 14354 36146 14366
rect 36206 14418 36258 14430
rect 36206 14354 36258 14366
rect 37102 14418 37154 14430
rect 37102 14354 37154 14366
rect 37662 14418 37714 14430
rect 45950 14418 46002 14430
rect 38882 14366 38894 14418
rect 38946 14366 38958 14418
rect 40786 14366 40798 14418
rect 40850 14366 40862 14418
rect 43138 14366 43150 14418
rect 43202 14366 43214 14418
rect 37662 14354 37714 14366
rect 45950 14354 46002 14366
rect 46734 14418 46786 14430
rect 46734 14354 46786 14366
rect 47966 14418 48018 14430
rect 47966 14354 48018 14366
rect 50878 14418 50930 14430
rect 50878 14354 50930 14366
rect 54574 14418 54626 14430
rect 54574 14354 54626 14366
rect 6974 14306 7026 14318
rect 6974 14242 7026 14254
rect 9886 14306 9938 14318
rect 26014 14306 26066 14318
rect 20178 14254 20190 14306
rect 20242 14254 20254 14306
rect 22754 14254 22766 14306
rect 22818 14254 22830 14306
rect 9886 14242 9938 14254
rect 26014 14242 26066 14254
rect 28030 14306 28082 14318
rect 28030 14242 28082 14254
rect 28254 14306 28306 14318
rect 28254 14242 28306 14254
rect 29150 14306 29202 14318
rect 29150 14242 29202 14254
rect 34974 14306 35026 14318
rect 34974 14242 35026 14254
rect 35422 14306 35474 14318
rect 35422 14242 35474 14254
rect 37886 14306 37938 14318
rect 37886 14242 37938 14254
rect 42814 14306 42866 14318
rect 42814 14242 42866 14254
rect 43486 14306 43538 14318
rect 43486 14242 43538 14254
rect 46510 14306 46562 14318
rect 46510 14242 46562 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 5966 13970 6018 13982
rect 5966 13906 6018 13918
rect 11566 13970 11618 13982
rect 24670 13970 24722 13982
rect 15474 13918 15486 13970
rect 15538 13918 15550 13970
rect 11566 13906 11618 13918
rect 24670 13906 24722 13918
rect 25678 13970 25730 13982
rect 25678 13906 25730 13918
rect 30270 13970 30322 13982
rect 43474 13918 43486 13970
rect 43538 13918 43550 13970
rect 30270 13906 30322 13918
rect 10222 13858 10274 13870
rect 10222 13794 10274 13806
rect 12014 13858 12066 13870
rect 18174 13858 18226 13870
rect 14466 13806 14478 13858
rect 14530 13806 14542 13858
rect 12014 13794 12066 13806
rect 18174 13794 18226 13806
rect 25454 13858 25506 13870
rect 25454 13794 25506 13806
rect 25902 13858 25954 13870
rect 25902 13794 25954 13806
rect 30830 13858 30882 13870
rect 46062 13858 46114 13870
rect 32498 13806 32510 13858
rect 32562 13806 32574 13858
rect 41794 13806 41806 13858
rect 41858 13806 41870 13858
rect 30830 13794 30882 13806
rect 46062 13794 46114 13806
rect 51774 13858 51826 13870
rect 51774 13794 51826 13806
rect 52222 13858 52274 13870
rect 52222 13794 52274 13806
rect 8430 13746 8482 13758
rect 13246 13746 13298 13758
rect 16830 13746 16882 13758
rect 7970 13694 7982 13746
rect 8034 13694 8046 13746
rect 9762 13694 9774 13746
rect 9826 13694 9838 13746
rect 10658 13694 10670 13746
rect 10722 13694 10734 13746
rect 11442 13694 11454 13746
rect 11506 13694 11518 13746
rect 14690 13694 14702 13746
rect 14754 13694 14766 13746
rect 15586 13694 15598 13746
rect 15650 13694 15662 13746
rect 8430 13682 8482 13694
rect 13246 13682 13298 13694
rect 16830 13682 16882 13694
rect 17838 13746 17890 13758
rect 20526 13746 20578 13758
rect 28366 13746 28418 13758
rect 38446 13746 38498 13758
rect 18050 13694 18062 13746
rect 18114 13694 18126 13746
rect 19506 13694 19518 13746
rect 19570 13694 19582 13746
rect 20962 13694 20974 13746
rect 21026 13694 21038 13746
rect 23314 13694 23326 13746
rect 23378 13694 23390 13746
rect 23538 13694 23550 13746
rect 23602 13694 23614 13746
rect 27682 13694 27694 13746
rect 27746 13694 27758 13746
rect 28914 13694 28926 13746
rect 28978 13694 28990 13746
rect 31042 13694 31054 13746
rect 31106 13694 31118 13746
rect 32162 13694 32174 13746
rect 32226 13694 32238 13746
rect 33730 13694 33742 13746
rect 33794 13694 33806 13746
rect 34738 13694 34750 13746
rect 34802 13694 34814 13746
rect 35522 13694 35534 13746
rect 35586 13694 35598 13746
rect 36978 13694 36990 13746
rect 37042 13694 37054 13746
rect 17838 13682 17890 13694
rect 20526 13682 20578 13694
rect 28366 13682 28418 13694
rect 38446 13682 38498 13694
rect 39902 13746 39954 13758
rect 39902 13682 39954 13694
rect 40014 13746 40066 13758
rect 43026 13694 43038 13746
rect 43090 13694 43102 13746
rect 45378 13694 45390 13746
rect 45442 13694 45454 13746
rect 51986 13694 51998 13746
rect 52050 13694 52062 13746
rect 40014 13682 40066 13694
rect 6526 13634 6578 13646
rect 6526 13570 6578 13582
rect 7086 13634 7138 13646
rect 7086 13570 7138 13582
rect 7534 13634 7586 13646
rect 7534 13570 7586 13582
rect 8990 13634 9042 13646
rect 8990 13570 9042 13582
rect 11118 13634 11170 13646
rect 11118 13570 11170 13582
rect 16270 13634 16322 13646
rect 16270 13570 16322 13582
rect 18734 13634 18786 13646
rect 33182 13634 33234 13646
rect 41022 13634 41074 13646
rect 21186 13582 21198 13634
rect 21250 13582 21262 13634
rect 23762 13582 23774 13634
rect 23826 13582 23838 13634
rect 25778 13582 25790 13634
rect 25842 13582 25854 13634
rect 27570 13582 27582 13634
rect 27634 13582 27646 13634
rect 31714 13582 31726 13634
rect 31778 13582 31790 13634
rect 37090 13582 37102 13634
rect 37154 13582 37166 13634
rect 38882 13582 38894 13634
rect 38946 13582 38958 13634
rect 18734 13570 18786 13582
rect 33182 13570 33234 13582
rect 41022 13570 41074 13582
rect 41694 13634 41746 13646
rect 45602 13582 45614 13634
rect 45666 13582 45678 13634
rect 51874 13582 51886 13634
rect 51938 13582 51950 13634
rect 41694 13570 41746 13582
rect 7198 13522 7250 13534
rect 20402 13470 20414 13522
rect 20466 13470 20478 13522
rect 23874 13470 23886 13522
rect 23938 13470 23950 13522
rect 29250 13470 29262 13522
rect 29314 13470 29326 13522
rect 37538 13470 37550 13522
rect 37602 13470 37614 13522
rect 38658 13470 38670 13522
rect 38722 13470 38734 13522
rect 7198 13458 7250 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 14030 13186 14082 13198
rect 18274 13134 18286 13186
rect 18338 13134 18350 13186
rect 32946 13134 32958 13186
rect 33010 13134 33022 13186
rect 14030 13122 14082 13134
rect 6750 13074 6802 13086
rect 6750 13010 6802 13022
rect 12910 13074 12962 13086
rect 12910 13010 12962 13022
rect 13806 13074 13858 13086
rect 35086 13074 35138 13086
rect 37550 13074 37602 13086
rect 41582 13074 41634 13086
rect 15810 13022 15822 13074
rect 15874 13022 15886 13074
rect 22642 13022 22654 13074
rect 22706 13022 22718 13074
rect 25106 13022 25118 13074
rect 25170 13022 25182 13074
rect 26226 13022 26238 13074
rect 26290 13022 26302 13074
rect 31938 13022 31950 13074
rect 32002 13022 32014 13074
rect 33730 13022 33742 13074
rect 33794 13022 33806 13074
rect 35858 13022 35870 13074
rect 35922 13022 35934 13074
rect 40898 13022 40910 13074
rect 40962 13022 40974 13074
rect 13806 13010 13858 13022
rect 35086 13010 35138 13022
rect 37550 13010 37602 13022
rect 41582 13010 41634 13022
rect 42366 13074 42418 13086
rect 57934 13074 57986 13086
rect 43362 13022 43374 13074
rect 43426 13022 43438 13074
rect 46946 13022 46958 13074
rect 47010 13022 47022 13074
rect 52770 13022 52782 13074
rect 52834 13022 52846 13074
rect 42366 13010 42418 13022
rect 57934 13010 57986 13022
rect 21870 12962 21922 12974
rect 26910 12962 26962 12974
rect 28030 12962 28082 12974
rect 6290 12910 6302 12962
rect 6354 12910 6366 12962
rect 7074 12910 7086 12962
rect 7138 12910 7150 12962
rect 8530 12910 8542 12962
rect 8594 12910 8606 12962
rect 10210 12910 10222 12962
rect 10274 12910 10286 12962
rect 12114 12910 12126 12962
rect 12178 12910 12190 12962
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 15026 12910 15038 12962
rect 15090 12910 15102 12962
rect 16930 12910 16942 12962
rect 16994 12910 17006 12962
rect 17602 12910 17614 12962
rect 17666 12910 17678 12962
rect 19058 12910 19070 12962
rect 19122 12910 19134 12962
rect 19842 12910 19854 12962
rect 19906 12910 19918 12962
rect 20626 12910 20638 12962
rect 20690 12910 20702 12962
rect 21410 12910 21422 12962
rect 21474 12910 21486 12962
rect 22978 12910 22990 12962
rect 23042 12910 23054 12962
rect 23986 12910 23998 12962
rect 24050 12910 24062 12962
rect 24994 12910 25006 12962
rect 25058 12910 25070 12962
rect 26114 12910 26126 12962
rect 26178 12910 26190 12962
rect 27346 12910 27358 12962
rect 27410 12910 27422 12962
rect 21870 12898 21922 12910
rect 26910 12898 26962 12910
rect 28030 12898 28082 12910
rect 28366 12962 28418 12974
rect 37886 12962 37938 12974
rect 44270 12962 44322 12974
rect 51326 12962 51378 12974
rect 28578 12910 28590 12962
rect 28642 12910 28654 12962
rect 29250 12910 29262 12962
rect 29314 12910 29326 12962
rect 30370 12910 30382 12962
rect 30434 12910 30446 12962
rect 31378 12910 31390 12962
rect 31442 12910 31454 12962
rect 32162 12910 32174 12962
rect 32226 12910 32238 12962
rect 32498 12910 32510 12962
rect 32562 12910 32574 12962
rect 33954 12910 33966 12962
rect 34018 12910 34030 12962
rect 34290 12910 34302 12962
rect 34354 12910 34366 12962
rect 38994 12910 39006 12962
rect 39058 12910 39070 12962
rect 39666 12910 39678 12962
rect 39730 12910 39742 12962
rect 40674 12910 40686 12962
rect 40738 12910 40750 12962
rect 43138 12910 43150 12962
rect 43202 12910 43214 12962
rect 46610 12910 46622 12962
rect 46674 12910 46686 12962
rect 28366 12898 28418 12910
rect 37886 12898 37938 12910
rect 44270 12898 44322 12910
rect 51326 12898 51378 12910
rect 51662 12962 51714 12974
rect 51662 12898 51714 12910
rect 51774 12962 51826 12974
rect 52994 12910 53006 12962
rect 53058 12910 53070 12962
rect 55906 12910 55918 12962
rect 55970 12910 55982 12962
rect 51774 12898 51826 12910
rect 22318 12850 22370 12862
rect 7410 12798 7422 12850
rect 7474 12798 7486 12850
rect 7858 12798 7870 12850
rect 7922 12798 7934 12850
rect 9650 12798 9662 12850
rect 9714 12798 9726 12850
rect 10098 12798 10110 12850
rect 10162 12798 10174 12850
rect 19730 12798 19742 12850
rect 19794 12798 19806 12850
rect 22318 12786 22370 12798
rect 22542 12850 22594 12862
rect 35534 12850 35586 12862
rect 24210 12798 24222 12850
rect 24274 12798 24286 12850
rect 24770 12798 24782 12850
rect 24834 12798 24846 12850
rect 26226 12798 26238 12850
rect 26290 12798 26302 12850
rect 33506 12798 33518 12850
rect 33570 12798 33582 12850
rect 22542 12786 22594 12798
rect 35534 12786 35586 12798
rect 37102 12850 37154 12862
rect 37102 12786 37154 12798
rect 38446 12850 38498 12862
rect 38446 12786 38498 12798
rect 41470 12850 41522 12862
rect 41470 12786 41522 12798
rect 41918 12850 41970 12862
rect 41918 12786 41970 12798
rect 43822 12850 43874 12862
rect 50990 12850 51042 12862
rect 49746 12798 49758 12850
rect 49810 12798 49822 12850
rect 43822 12786 43874 12798
rect 50990 12786 51042 12798
rect 51102 12850 51154 12862
rect 51102 12786 51154 12798
rect 52110 12850 52162 12862
rect 52110 12786 52162 12798
rect 53678 12850 53730 12862
rect 53678 12786 53730 12798
rect 12350 12738 12402 12750
rect 28142 12738 28194 12750
rect 8082 12686 8094 12738
rect 8146 12686 8158 12738
rect 20626 12686 20638 12738
rect 20690 12686 20702 12738
rect 12350 12674 12402 12686
rect 28142 12674 28194 12686
rect 28254 12738 28306 12750
rect 28254 12674 28306 12686
rect 31390 12738 31442 12750
rect 31390 12674 31442 12686
rect 35758 12738 35810 12750
rect 35758 12674 35810 12686
rect 36318 12738 36370 12750
rect 36318 12674 36370 12686
rect 38222 12738 38274 12750
rect 38222 12674 38274 12686
rect 38558 12738 38610 12750
rect 38558 12674 38610 12686
rect 41694 12738 41746 12750
rect 41694 12674 41746 12686
rect 49422 12738 49474 12750
rect 49422 12674 49474 12686
rect 51998 12738 52050 12750
rect 51998 12674 52050 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 9102 12402 9154 12414
rect 9102 12338 9154 12350
rect 9886 12402 9938 12414
rect 9886 12338 9938 12350
rect 37774 12402 37826 12414
rect 37774 12338 37826 12350
rect 38446 12402 38498 12414
rect 38446 12338 38498 12350
rect 39342 12402 39394 12414
rect 39342 12338 39394 12350
rect 39454 12402 39506 12414
rect 39454 12338 39506 12350
rect 40126 12402 40178 12414
rect 40126 12338 40178 12350
rect 42030 12402 42082 12414
rect 51886 12402 51938 12414
rect 50418 12350 50430 12402
rect 50482 12350 50494 12402
rect 42030 12338 42082 12350
rect 51886 12338 51938 12350
rect 52334 12402 52386 12414
rect 52334 12338 52386 12350
rect 55918 12402 55970 12414
rect 55918 12338 55970 12350
rect 16270 12290 16322 12302
rect 33070 12290 33122 12302
rect 7298 12238 7310 12290
rect 7362 12238 7374 12290
rect 10994 12238 11006 12290
rect 11058 12238 11070 12290
rect 12450 12238 12462 12290
rect 12514 12238 12526 12290
rect 13682 12238 13694 12290
rect 13746 12238 13758 12290
rect 26002 12238 26014 12290
rect 26066 12238 26078 12290
rect 30370 12238 30382 12290
rect 30434 12238 30446 12290
rect 16270 12226 16322 12238
rect 33070 12226 33122 12238
rect 34078 12290 34130 12302
rect 34078 12226 34130 12238
rect 35646 12290 35698 12302
rect 35646 12226 35698 12238
rect 37326 12290 37378 12302
rect 37326 12226 37378 12238
rect 40014 12290 40066 12302
rect 43934 12290 43986 12302
rect 41234 12238 41246 12290
rect 41298 12238 41310 12290
rect 40014 12226 40066 12238
rect 43934 12226 43986 12238
rect 46174 12290 46226 12302
rect 49982 12290 50034 12302
rect 52670 12290 52722 12302
rect 48178 12238 48190 12290
rect 48242 12238 48254 12290
rect 49074 12238 49086 12290
rect 49138 12238 49150 12290
rect 49298 12238 49310 12290
rect 49362 12238 49374 12290
rect 51090 12238 51102 12290
rect 51154 12238 51166 12290
rect 46174 12226 46226 12238
rect 49982 12226 50034 12238
rect 52670 12226 52722 12238
rect 53006 12290 53058 12302
rect 53006 12226 53058 12238
rect 6302 12178 6354 12190
rect 7982 12178 8034 12190
rect 22766 12178 22818 12190
rect 27134 12178 27186 12190
rect 35086 12178 35138 12190
rect 37550 12178 37602 12190
rect 5842 12126 5854 12178
rect 5906 12126 5918 12178
rect 7522 12126 7534 12178
rect 7586 12126 7598 12178
rect 10322 12126 10334 12178
rect 10386 12126 10398 12178
rect 10882 12126 10894 12178
rect 10946 12126 10958 12178
rect 11554 12126 11566 12178
rect 11618 12126 11630 12178
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 13234 12126 13246 12178
rect 13298 12126 13310 12178
rect 13570 12126 13582 12178
rect 13634 12126 13646 12178
rect 14578 12126 14590 12178
rect 14642 12126 14654 12178
rect 14802 12126 14814 12178
rect 14866 12126 14878 12178
rect 15922 12126 15934 12178
rect 15986 12126 15998 12178
rect 16706 12126 16718 12178
rect 16770 12126 16782 12178
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 19842 12126 19854 12178
rect 19906 12126 19918 12178
rect 20738 12126 20750 12178
rect 20802 12126 20814 12178
rect 21186 12126 21198 12178
rect 21250 12126 21262 12178
rect 24546 12126 24558 12178
rect 24610 12126 24622 12178
rect 26226 12126 26238 12178
rect 26290 12126 26302 12178
rect 27346 12126 27358 12178
rect 27410 12126 27422 12178
rect 29474 12126 29486 12178
rect 29538 12126 29550 12178
rect 29810 12126 29822 12178
rect 29874 12126 29886 12178
rect 30706 12126 30718 12178
rect 30770 12126 30782 12178
rect 31602 12126 31614 12178
rect 31666 12126 31678 12178
rect 33282 12126 33294 12178
rect 33346 12126 33358 12178
rect 34514 12126 34526 12178
rect 34578 12126 34590 12178
rect 36418 12126 36430 12178
rect 36482 12126 36494 12178
rect 6302 12114 6354 12126
rect 7982 12114 8034 12126
rect 22766 12114 22818 12126
rect 27134 12114 27186 12126
rect 35086 12114 35138 12126
rect 37550 12114 37602 12126
rect 37886 12178 37938 12190
rect 37886 12114 37938 12126
rect 38894 12178 38946 12190
rect 38894 12114 38946 12126
rect 39566 12178 39618 12190
rect 39566 12114 39618 12126
rect 42926 12178 42978 12190
rect 45390 12178 45442 12190
rect 52110 12178 52162 12190
rect 45042 12126 45054 12178
rect 45106 12126 45118 12178
rect 45714 12126 45726 12178
rect 45778 12126 45790 12178
rect 46946 12126 46958 12178
rect 47010 12126 47022 12178
rect 47506 12126 47518 12178
rect 47570 12126 47582 12178
rect 48850 12126 48862 12178
rect 48914 12126 48926 12178
rect 50194 12126 50206 12178
rect 50258 12126 50270 12178
rect 50754 12126 50766 12178
rect 50818 12126 50830 12178
rect 42926 12114 42978 12126
rect 45390 12114 45442 12126
rect 52110 12114 52162 12126
rect 52782 12178 52834 12190
rect 52782 12114 52834 12126
rect 53454 12178 53506 12190
rect 55246 12178 55298 12190
rect 54562 12126 54574 12178
rect 54626 12126 54638 12178
rect 53454 12114 53506 12126
rect 55246 12114 55298 12126
rect 55582 12178 55634 12190
rect 55582 12114 55634 12126
rect 6862 12066 6914 12078
rect 17726 12066 17778 12078
rect 52222 12066 52274 12078
rect 11106 12014 11118 12066
rect 11170 12014 11182 12066
rect 12562 12014 12574 12066
rect 12626 12014 12638 12066
rect 14018 12014 14030 12066
rect 14082 12014 14094 12066
rect 18610 12014 18622 12066
rect 18674 12014 18686 12066
rect 19730 12014 19742 12066
rect 19794 12014 19806 12066
rect 23202 12014 23214 12066
rect 23266 12014 23278 12066
rect 29698 12014 29710 12066
rect 29762 12014 29774 12066
rect 31378 12014 31390 12066
rect 31442 12014 31454 12066
rect 36866 12014 36878 12066
rect 36930 12014 36942 12066
rect 47394 12014 47406 12066
rect 47458 12014 47470 12066
rect 54338 12014 54350 12066
rect 54402 12014 54414 12066
rect 6862 12002 6914 12014
rect 17726 12002 17778 12014
rect 52222 12002 52274 12014
rect 8318 11954 8370 11966
rect 24446 11954 24498 11966
rect 40126 11954 40178 11966
rect 14802 11902 14814 11954
rect 14866 11902 14878 11954
rect 17378 11902 17390 11954
rect 17442 11951 17454 11954
rect 17714 11951 17726 11954
rect 17442 11905 17726 11951
rect 17442 11902 17454 11905
rect 17714 11902 17726 11905
rect 17778 11902 17790 11954
rect 23314 11902 23326 11954
rect 23378 11902 23390 11954
rect 28354 11902 28366 11954
rect 28418 11902 28430 11954
rect 31826 11902 31838 11954
rect 31890 11902 31902 11954
rect 33394 11902 33406 11954
rect 33458 11902 33470 11954
rect 8318 11890 8370 11902
rect 24446 11890 24498 11902
rect 40126 11890 40178 11902
rect 53230 11954 53282 11966
rect 53230 11890 53282 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 20078 11618 20130 11630
rect 30830 11618 30882 11630
rect 42814 11618 42866 11630
rect 9762 11615 9774 11618
rect 8657 11569 9774 11615
rect 7534 11506 7586 11518
rect 7534 11442 7586 11454
rect 8430 11506 8482 11518
rect 8657 11506 8703 11569
rect 9762 11566 9774 11569
rect 9826 11566 9838 11618
rect 10658 11615 10670 11618
rect 10337 11569 10670 11615
rect 8766 11506 8818 11518
rect 8642 11454 8654 11506
rect 8706 11454 8718 11506
rect 8430 11442 8482 11454
rect 8766 11442 8818 11454
rect 10110 11506 10162 11518
rect 10337 11506 10383 11569
rect 10658 11566 10670 11569
rect 10722 11566 10734 11618
rect 25106 11566 25118 11618
rect 25170 11566 25182 11618
rect 39666 11615 39678 11618
rect 20078 11554 20130 11566
rect 30830 11554 30882 11566
rect 39233 11569 39678 11615
rect 12574 11506 12626 11518
rect 19070 11506 19122 11518
rect 10322 11454 10334 11506
rect 10386 11454 10398 11506
rect 14018 11454 14030 11506
rect 14082 11454 14094 11506
rect 10110 11442 10162 11454
rect 12574 11442 12626 11454
rect 19070 11442 19122 11454
rect 21870 11506 21922 11518
rect 31390 11506 31442 11518
rect 24434 11454 24446 11506
rect 24498 11454 24510 11506
rect 27122 11454 27134 11506
rect 27186 11454 27198 11506
rect 21870 11442 21922 11454
rect 31390 11442 31442 11454
rect 38446 11506 38498 11518
rect 38882 11454 38894 11506
rect 38946 11503 38958 11506
rect 39233 11503 39279 11569
rect 39666 11566 39678 11569
rect 39730 11615 39742 11618
rect 40226 11615 40238 11618
rect 39730 11569 40238 11615
rect 39730 11566 39742 11569
rect 40226 11566 40238 11569
rect 40290 11566 40302 11618
rect 40450 11566 40462 11618
rect 40514 11615 40526 11618
rect 41234 11615 41246 11618
rect 40514 11569 41246 11615
rect 40514 11566 40526 11569
rect 41234 11566 41246 11569
rect 41298 11566 41310 11618
rect 42814 11554 42866 11566
rect 47182 11618 47234 11630
rect 47182 11554 47234 11566
rect 48302 11618 48354 11630
rect 48302 11554 48354 11566
rect 54350 11618 54402 11630
rect 54350 11554 54402 11566
rect 38946 11457 39279 11503
rect 39902 11506 39954 11518
rect 38946 11454 38958 11457
rect 38446 11442 38498 11454
rect 39902 11442 39954 11454
rect 40238 11506 40290 11518
rect 40238 11442 40290 11454
rect 41246 11506 41298 11518
rect 46398 11506 46450 11518
rect 43586 11454 43598 11506
rect 43650 11454 43662 11506
rect 41246 11442 41298 11454
rect 46398 11442 46450 11454
rect 46734 11506 46786 11518
rect 53902 11506 53954 11518
rect 52994 11454 53006 11506
rect 53058 11454 53070 11506
rect 46734 11442 46786 11454
rect 53902 11442 53954 11454
rect 21310 11394 21362 11406
rect 29486 11394 29538 11406
rect 31726 11394 31778 11406
rect 37102 11394 37154 11406
rect 37998 11394 38050 11406
rect 11106 11342 11118 11394
rect 11170 11342 11182 11394
rect 11554 11342 11566 11394
rect 11618 11342 11630 11394
rect 12114 11342 12126 11394
rect 12178 11342 12190 11394
rect 13682 11342 13694 11394
rect 13746 11342 13758 11394
rect 14914 11342 14926 11394
rect 14978 11342 14990 11394
rect 16258 11342 16270 11394
rect 16322 11342 16334 11394
rect 16818 11342 16830 11394
rect 16882 11342 16894 11394
rect 19170 11342 19182 11394
rect 19234 11342 19246 11394
rect 19954 11342 19966 11394
rect 20018 11342 20030 11394
rect 23426 11342 23438 11394
rect 23490 11342 23502 11394
rect 24322 11342 24334 11394
rect 24386 11342 24398 11394
rect 26114 11342 26126 11394
rect 26178 11342 26190 11394
rect 27234 11342 27246 11394
rect 27298 11342 27310 11394
rect 27794 11342 27806 11394
rect 27858 11342 27870 11394
rect 28242 11342 28254 11394
rect 28306 11342 28318 11394
rect 30818 11342 30830 11394
rect 30882 11342 30894 11394
rect 32386 11342 32398 11394
rect 32450 11342 32462 11394
rect 34626 11342 34638 11394
rect 34690 11342 34702 11394
rect 36306 11342 36318 11394
rect 36370 11342 36382 11394
rect 37538 11342 37550 11394
rect 37602 11342 37614 11394
rect 21310 11330 21362 11342
rect 29486 11330 29538 11342
rect 31726 11330 31778 11342
rect 37102 11330 37154 11342
rect 37998 11330 38050 11342
rect 42030 11394 42082 11406
rect 42030 11330 42082 11342
rect 42254 11394 42306 11406
rect 46958 11394 47010 11406
rect 43362 11342 43374 11394
rect 43426 11342 43438 11394
rect 42254 11330 42306 11342
rect 46958 11330 47010 11342
rect 47630 11394 47682 11406
rect 47630 11330 47682 11342
rect 47966 11394 48018 11406
rect 47966 11330 48018 11342
rect 48190 11394 48242 11406
rect 49310 11394 49362 11406
rect 49074 11342 49086 11394
rect 49138 11342 49150 11394
rect 48190 11330 48242 11342
rect 49310 11330 49362 11342
rect 49422 11394 49474 11406
rect 49422 11330 49474 11342
rect 54238 11394 54290 11406
rect 54238 11330 54290 11342
rect 10670 11282 10722 11294
rect 10670 11218 10722 11230
rect 11678 11282 11730 11294
rect 28366 11282 28418 11294
rect 17602 11230 17614 11282
rect 17666 11230 17678 11282
rect 22978 11230 22990 11282
rect 23042 11230 23054 11282
rect 27010 11230 27022 11282
rect 27074 11230 27086 11282
rect 11678 11218 11730 11230
rect 28366 11218 28418 11230
rect 29262 11282 29314 11294
rect 29262 11218 29314 11230
rect 29374 11282 29426 11294
rect 29374 11218 29426 11230
rect 30494 11282 30546 11294
rect 30494 11218 30546 11230
rect 32062 11282 32114 11294
rect 38782 11282 38834 11294
rect 32274 11230 32286 11282
rect 32338 11230 32350 11282
rect 36418 11230 36430 11282
rect 36482 11230 36494 11282
rect 32062 11218 32114 11230
rect 38782 11218 38834 11230
rect 42590 11282 42642 11294
rect 42590 11218 42642 11230
rect 44270 11282 44322 11294
rect 44270 11218 44322 11230
rect 47854 11282 47906 11294
rect 52770 11230 52782 11282
rect 52834 11230 52846 11282
rect 47854 11218 47906 11230
rect 6638 11170 6690 11182
rect 6638 11106 6690 11118
rect 6974 11170 7026 11182
rect 6974 11106 7026 11118
rect 7982 11170 8034 11182
rect 7982 11106 8034 11118
rect 9326 11170 9378 11182
rect 9326 11106 9378 11118
rect 9662 11170 9714 11182
rect 9662 11106 9714 11118
rect 18062 11170 18114 11182
rect 18062 11106 18114 11118
rect 20750 11170 20802 11182
rect 31838 11170 31890 11182
rect 38334 11170 38386 11182
rect 29922 11118 29934 11170
rect 29986 11118 29998 11170
rect 36194 11118 36206 11170
rect 36258 11118 36270 11170
rect 20750 11106 20802 11118
rect 31838 11106 31890 11118
rect 38334 11106 38386 11118
rect 38558 11170 38610 11182
rect 38558 11106 38610 11118
rect 39342 11170 39394 11182
rect 39342 11106 39394 11118
rect 40686 11170 40738 11182
rect 40686 11106 40738 11118
rect 41918 11170 41970 11182
rect 49858 11118 49870 11170
rect 49922 11118 49934 11170
rect 41918 11106 41970 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 7086 10834 7138 10846
rect 7086 10770 7138 10782
rect 8094 10834 8146 10846
rect 8094 10770 8146 10782
rect 10110 10834 10162 10846
rect 14478 10834 14530 10846
rect 13906 10782 13918 10834
rect 13970 10782 13982 10834
rect 10110 10770 10162 10782
rect 14478 10770 14530 10782
rect 17726 10834 17778 10846
rect 24110 10834 24162 10846
rect 21634 10782 21646 10834
rect 21698 10782 21710 10834
rect 17726 10770 17778 10782
rect 24110 10770 24162 10782
rect 24222 10834 24274 10846
rect 24222 10770 24274 10782
rect 27582 10834 27634 10846
rect 35086 10834 35138 10846
rect 41694 10834 41746 10846
rect 32386 10782 32398 10834
rect 32450 10782 32462 10834
rect 37202 10782 37214 10834
rect 37266 10782 37278 10834
rect 27582 10770 27634 10782
rect 35086 10770 35138 10782
rect 41694 10770 41746 10782
rect 42814 10834 42866 10846
rect 42814 10770 42866 10782
rect 43374 10834 43426 10846
rect 43374 10770 43426 10782
rect 43598 10834 43650 10846
rect 43598 10770 43650 10782
rect 45950 10834 46002 10846
rect 45950 10770 46002 10782
rect 50094 10834 50146 10846
rect 50094 10770 50146 10782
rect 50318 10834 50370 10846
rect 50318 10770 50370 10782
rect 51998 10834 52050 10846
rect 51998 10770 52050 10782
rect 53790 10834 53842 10846
rect 53790 10770 53842 10782
rect 8542 10722 8594 10734
rect 12910 10722 12962 10734
rect 25230 10722 25282 10734
rect 36206 10722 36258 10734
rect 10322 10670 10334 10722
rect 10386 10670 10398 10722
rect 20850 10670 20862 10722
rect 20914 10670 20926 10722
rect 22978 10670 22990 10722
rect 23042 10670 23054 10722
rect 26002 10670 26014 10722
rect 26066 10670 26078 10722
rect 28578 10670 28590 10722
rect 28642 10670 28654 10722
rect 31602 10670 31614 10722
rect 31666 10670 31678 10722
rect 34514 10670 34526 10722
rect 34578 10670 34590 10722
rect 8542 10658 8594 10670
rect 12910 10658 12962 10670
rect 25230 10658 25282 10670
rect 36206 10658 36258 10670
rect 38222 10722 38274 10734
rect 53006 10722 53058 10734
rect 48178 10670 48190 10722
rect 48242 10670 48254 10722
rect 38222 10658 38274 10670
rect 53006 10658 53058 10670
rect 53566 10722 53618 10734
rect 53566 10658 53618 10670
rect 6526 10610 6578 10622
rect 7758 10610 7810 10622
rect 5730 10558 5742 10610
rect 5794 10558 5806 10610
rect 7522 10558 7534 10610
rect 7586 10558 7598 10610
rect 6526 10546 6578 10558
rect 7758 10546 7810 10558
rect 12014 10610 12066 10622
rect 15262 10610 15314 10622
rect 12338 10558 12350 10610
rect 12402 10558 12414 10610
rect 12014 10546 12066 10558
rect 15262 10546 15314 10558
rect 15598 10610 15650 10622
rect 15598 10546 15650 10558
rect 15822 10610 15874 10622
rect 17950 10610 18002 10622
rect 16706 10558 16718 10610
rect 16770 10558 16782 10610
rect 15822 10546 15874 10558
rect 17950 10546 18002 10558
rect 18174 10610 18226 10622
rect 24334 10610 24386 10622
rect 26238 10610 26290 10622
rect 43262 10610 43314 10622
rect 18610 10558 18622 10610
rect 18674 10558 18686 10610
rect 19170 10558 19182 10610
rect 19234 10558 19246 10610
rect 19730 10558 19742 10610
rect 19794 10558 19806 10610
rect 20962 10558 20974 10610
rect 21026 10558 21038 10610
rect 22194 10558 22206 10610
rect 22258 10558 22270 10610
rect 24658 10558 24670 10610
rect 24722 10558 24734 10610
rect 25442 10558 25454 10610
rect 25506 10558 25518 10610
rect 26674 10558 26686 10610
rect 26738 10558 26750 10610
rect 28802 10558 28814 10610
rect 28866 10558 28878 10610
rect 29810 10558 29822 10610
rect 29874 10558 29886 10610
rect 30258 10558 30270 10610
rect 30322 10558 30334 10610
rect 31378 10558 31390 10610
rect 31442 10558 31454 10610
rect 32274 10558 32286 10610
rect 32338 10558 32350 10610
rect 33394 10558 33406 10610
rect 33458 10558 33470 10610
rect 34290 10558 34302 10610
rect 34354 10558 34366 10610
rect 35634 10558 35646 10610
rect 35698 10558 35710 10610
rect 37650 10558 37662 10610
rect 37714 10558 37726 10610
rect 41234 10558 41246 10610
rect 41298 10558 41310 10610
rect 18174 10546 18226 10558
rect 24334 10546 24386 10558
rect 26238 10546 26290 10558
rect 43262 10546 43314 10558
rect 44830 10610 44882 10622
rect 49646 10610 49698 10622
rect 45154 10558 45166 10610
rect 45218 10558 45230 10610
rect 46722 10558 46734 10610
rect 46786 10558 46798 10610
rect 47506 10558 47518 10610
rect 47570 10558 47582 10610
rect 48066 10558 48078 10610
rect 48130 10558 48142 10610
rect 44830 10546 44882 10558
rect 49646 10546 49698 10558
rect 51102 10610 51154 10622
rect 51202 10558 51214 10610
rect 51266 10558 51278 10610
rect 51102 10546 51154 10558
rect 6190 10498 6242 10510
rect 6190 10434 6242 10446
rect 15038 10498 15090 10510
rect 15038 10434 15090 10446
rect 15486 10498 15538 10510
rect 15486 10434 15538 10446
rect 16270 10498 16322 10510
rect 16270 10434 16322 10446
rect 18062 10498 18114 10510
rect 18062 10434 18114 10446
rect 28142 10498 28194 10510
rect 28142 10434 28194 10446
rect 28702 10498 28754 10510
rect 28702 10434 28754 10446
rect 30718 10498 30770 10510
rect 50206 10498 50258 10510
rect 52782 10498 52834 10510
rect 33842 10446 33854 10498
rect 33906 10446 33918 10498
rect 42914 10446 42926 10498
rect 42978 10446 42990 10498
rect 46386 10446 46398 10498
rect 46450 10446 46462 10498
rect 50754 10446 50766 10498
rect 50818 10446 50830 10498
rect 53106 10446 53118 10498
rect 53170 10446 53182 10498
rect 53890 10446 53902 10498
rect 53954 10446 53966 10498
rect 30718 10434 30770 10446
rect 50206 10434 50258 10446
rect 52782 10434 52834 10446
rect 8654 10386 8706 10398
rect 8654 10322 8706 10334
rect 19406 10386 19458 10398
rect 19406 10322 19458 10334
rect 40910 10386 40962 10398
rect 40910 10322 40962 10334
rect 41246 10386 41298 10398
rect 41246 10322 41298 10334
rect 42590 10386 42642 10398
rect 45490 10334 45502 10386
rect 45554 10334 45566 10386
rect 42590 10322 42642 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 13694 10050 13746 10062
rect 28366 10050 28418 10062
rect 46846 10050 46898 10062
rect 16146 9998 16158 10050
rect 16210 9998 16222 10050
rect 20402 9998 20414 10050
rect 20466 9998 20478 10050
rect 22194 9998 22206 10050
rect 22258 9998 22270 10050
rect 27346 9998 27358 10050
rect 27410 9998 27422 10050
rect 33394 9998 33406 10050
rect 33458 9998 33470 10050
rect 13694 9986 13746 9998
rect 28366 9986 28418 9998
rect 46846 9986 46898 9998
rect 47070 10050 47122 10062
rect 47070 9986 47122 9998
rect 50766 10050 50818 10062
rect 50766 9986 50818 9998
rect 50990 10050 51042 10062
rect 50990 9986 51042 9998
rect 5966 9938 6018 9950
rect 24670 9938 24722 9950
rect 35758 9938 35810 9950
rect 38558 9938 38610 9950
rect 7858 9886 7870 9938
rect 7922 9886 7934 9938
rect 9874 9886 9886 9938
rect 9938 9886 9950 9938
rect 14690 9886 14702 9938
rect 14754 9886 14766 9938
rect 20178 9886 20190 9938
rect 20242 9886 20254 9938
rect 23090 9886 23102 9938
rect 23154 9886 23166 9938
rect 32946 9886 32958 9938
rect 33010 9886 33022 9938
rect 34738 9886 34750 9938
rect 34802 9886 34814 9938
rect 37090 9886 37102 9938
rect 37154 9886 37166 9938
rect 5966 9874 6018 9886
rect 24670 9874 24722 9886
rect 35758 9874 35810 9886
rect 38558 9874 38610 9886
rect 41470 9938 41522 9950
rect 41470 9874 41522 9886
rect 45838 9938 45890 9950
rect 50542 9938 50594 9950
rect 48626 9886 48638 9938
rect 48690 9886 48702 9938
rect 45838 9874 45890 9886
rect 50542 9874 50594 9886
rect 51438 9938 51490 9950
rect 51438 9874 51490 9886
rect 12238 9826 12290 9838
rect 7746 9774 7758 9826
rect 7810 9774 7822 9826
rect 9426 9774 9438 9826
rect 9490 9774 9502 9826
rect 10546 9774 10558 9826
rect 10610 9774 10622 9826
rect 12238 9762 12290 9774
rect 12910 9826 12962 9838
rect 12910 9762 12962 9774
rect 13806 9826 13858 9838
rect 22094 9826 22146 9838
rect 14354 9774 14366 9826
rect 14418 9774 14430 9826
rect 16034 9774 16046 9826
rect 16098 9774 16110 9826
rect 17378 9774 17390 9826
rect 17442 9774 17454 9826
rect 18498 9774 18510 9826
rect 18562 9774 18574 9826
rect 19618 9774 19630 9826
rect 19682 9774 19694 9826
rect 20402 9774 20414 9826
rect 20466 9774 20478 9826
rect 21746 9774 21758 9826
rect 21810 9774 21822 9826
rect 13806 9762 13858 9774
rect 22094 9762 22146 9774
rect 22654 9826 22706 9838
rect 22654 9762 22706 9774
rect 23886 9826 23938 9838
rect 26238 9826 26290 9838
rect 24210 9774 24222 9826
rect 24274 9774 24286 9826
rect 25106 9774 25118 9826
rect 25170 9774 25182 9826
rect 23886 9762 23938 9774
rect 26238 9762 26290 9774
rect 26686 9826 26738 9838
rect 28030 9826 28082 9838
rect 27010 9774 27022 9826
rect 27074 9774 27086 9826
rect 27794 9774 27806 9826
rect 27858 9774 27870 9826
rect 26686 9762 26738 9774
rect 28030 9762 28082 9774
rect 28254 9826 28306 9838
rect 34302 9826 34354 9838
rect 37998 9826 38050 9838
rect 29586 9774 29598 9826
rect 29650 9774 29662 9826
rect 29922 9774 29934 9826
rect 29986 9774 29998 9826
rect 31378 9774 31390 9826
rect 31442 9774 31454 9826
rect 32498 9774 32510 9826
rect 32562 9774 32574 9826
rect 37426 9774 37438 9826
rect 37490 9774 37502 9826
rect 28254 9762 28306 9774
rect 34302 9762 34354 9774
rect 37998 9762 38050 9774
rect 39566 9826 39618 9838
rect 39566 9762 39618 9774
rect 39902 9826 39954 9838
rect 46622 9826 46674 9838
rect 40338 9774 40350 9826
rect 40402 9774 40414 9826
rect 41794 9774 41806 9826
rect 41858 9774 41870 9826
rect 42242 9774 42254 9826
rect 42306 9774 42318 9826
rect 47842 9774 47854 9826
rect 47906 9774 47918 9826
rect 48402 9774 48414 9826
rect 48466 9774 48478 9826
rect 39902 9762 39954 9774
rect 46622 9762 46674 9774
rect 12686 9714 12738 9726
rect 11666 9662 11678 9714
rect 11730 9662 11742 9714
rect 12686 9650 12738 9662
rect 17166 9714 17218 9726
rect 18174 9714 18226 9726
rect 17714 9662 17726 9714
rect 17778 9662 17790 9714
rect 17166 9650 17218 9662
rect 18174 9650 18226 9662
rect 39342 9714 39394 9726
rect 41694 9714 41746 9726
rect 40562 9662 40574 9714
rect 40626 9662 40638 9714
rect 41010 9662 41022 9714
rect 41074 9662 41086 9714
rect 39342 9650 39394 9662
rect 41694 9650 41746 9662
rect 42814 9714 42866 9726
rect 51662 9714 51714 9726
rect 48962 9662 48974 9714
rect 49026 9662 49038 9714
rect 42814 9650 42866 9662
rect 51662 9650 51714 9662
rect 51774 9714 51826 9726
rect 51774 9650 51826 9662
rect 6414 9602 6466 9614
rect 6414 9538 6466 9550
rect 6862 9602 6914 9614
rect 6862 9538 6914 9550
rect 7310 9602 7362 9614
rect 7310 9538 7362 9550
rect 12798 9602 12850 9614
rect 12798 9538 12850 9550
rect 13694 9602 13746 9614
rect 13694 9538 13746 9550
rect 35310 9602 35362 9614
rect 35310 9538 35362 9550
rect 36206 9602 36258 9614
rect 36206 9538 36258 9550
rect 39566 9602 39618 9614
rect 39566 9538 39618 9550
rect 42926 9602 42978 9614
rect 42926 9538 42978 9550
rect 43150 9602 43202 9614
rect 43150 9538 43202 9550
rect 43486 9602 43538 9614
rect 43486 9538 43538 9550
rect 47518 9602 47570 9614
rect 47518 9538 47570 9550
rect 51998 9602 52050 9614
rect 51998 9538 52050 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 6526 9266 6578 9278
rect 6526 9202 6578 9214
rect 6862 9266 6914 9278
rect 6862 9202 6914 9214
rect 9102 9266 9154 9278
rect 9102 9202 9154 9214
rect 9550 9266 9602 9278
rect 9550 9202 9602 9214
rect 10446 9266 10498 9278
rect 17614 9266 17666 9278
rect 14914 9214 14926 9266
rect 14978 9214 14990 9266
rect 10446 9202 10498 9214
rect 17614 9202 17666 9214
rect 22654 9266 22706 9278
rect 22654 9202 22706 9214
rect 22766 9266 22818 9278
rect 27694 9266 27746 9278
rect 24098 9214 24110 9266
rect 24162 9214 24174 9266
rect 22766 9202 22818 9214
rect 27694 9202 27746 9214
rect 29598 9266 29650 9278
rect 39118 9266 39170 9278
rect 34066 9214 34078 9266
rect 34130 9214 34142 9266
rect 29598 9202 29650 9214
rect 39118 9202 39170 9214
rect 39566 9266 39618 9278
rect 39566 9202 39618 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 44158 9266 44210 9278
rect 44158 9202 44210 9214
rect 45614 9266 45666 9278
rect 45614 9202 45666 9214
rect 1710 9154 1762 9166
rect 10222 9154 10274 9166
rect 17838 9154 17890 9166
rect 42030 9154 42082 9166
rect 7858 9102 7870 9154
rect 7922 9102 7934 9154
rect 8306 9102 8318 9154
rect 8370 9102 8382 9154
rect 9874 9102 9886 9154
rect 9938 9102 9950 9154
rect 13682 9102 13694 9154
rect 13746 9102 13758 9154
rect 14130 9102 14142 9154
rect 14194 9102 14206 9154
rect 20738 9102 20750 9154
rect 20802 9102 20814 9154
rect 23314 9102 23326 9154
rect 23378 9102 23390 9154
rect 25554 9102 25566 9154
rect 25618 9102 25630 9154
rect 28018 9102 28030 9154
rect 28082 9102 28094 9154
rect 31490 9102 31502 9154
rect 31554 9102 31566 9154
rect 33170 9102 33182 9154
rect 33234 9102 33246 9154
rect 35858 9102 35870 9154
rect 35922 9102 35934 9154
rect 36978 9102 36990 9154
rect 37042 9102 37054 9154
rect 38770 9102 38782 9154
rect 38834 9102 38846 9154
rect 1710 9090 1762 9102
rect 10222 9090 10274 9102
rect 17838 9090 17890 9102
rect 42030 9090 42082 9102
rect 44606 9154 44658 9166
rect 44606 9090 44658 9102
rect 44830 9154 44882 9166
rect 44830 9090 44882 9102
rect 48750 9154 48802 9166
rect 48750 9090 48802 9102
rect 48862 9154 48914 9166
rect 48862 9090 48914 9102
rect 54014 9154 54066 9166
rect 54014 9090 54066 9102
rect 6190 9042 6242 9054
rect 27134 9042 27186 9054
rect 49086 9042 49138 9054
rect 53342 9042 53394 9054
rect 7746 8990 7758 9042
rect 7810 8990 7822 9042
rect 11218 8990 11230 9042
rect 11282 8990 11294 9042
rect 11890 8990 11902 9042
rect 11954 8990 11966 9042
rect 12562 8990 12574 9042
rect 12626 8990 12638 9042
rect 13122 8990 13134 9042
rect 13186 8990 13198 9042
rect 14578 8990 14590 9042
rect 14642 8990 14654 9042
rect 14914 8990 14926 9042
rect 14978 8990 14990 9042
rect 15922 8990 15934 9042
rect 15986 8990 15998 9042
rect 16258 8990 16270 9042
rect 16322 8990 16334 9042
rect 19506 8990 19518 9042
rect 19570 8990 19582 9042
rect 21074 8990 21086 9042
rect 21138 8990 21150 9042
rect 21858 8990 21870 9042
rect 21922 8990 21934 9042
rect 23650 8990 23662 9042
rect 23714 8990 23726 9042
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 25442 8990 25454 9042
rect 25506 8990 25518 9042
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 29810 8990 29822 9042
rect 29874 8990 29886 9042
rect 31826 8990 31838 9042
rect 31890 8990 31902 9042
rect 33058 8990 33070 9042
rect 33122 8990 33134 9042
rect 34178 8990 34190 9042
rect 34242 8990 34254 9042
rect 36306 8990 36318 9042
rect 36370 8990 36382 9042
rect 36754 8990 36766 9042
rect 36818 8990 36830 9042
rect 41234 8990 41246 9042
rect 41298 8990 41310 9042
rect 52658 8990 52670 9042
rect 52722 8990 52734 9042
rect 6190 8978 6242 8990
rect 27134 8978 27186 8990
rect 49086 8978 49138 8990
rect 53342 8978 53394 8990
rect 53678 9042 53730 9054
rect 53678 8978 53730 8990
rect 7422 8930 7474 8942
rect 20526 8930 20578 8942
rect 34638 8930 34690 8942
rect 42814 8930 42866 8942
rect 10994 8878 11006 8930
rect 11058 8878 11070 8930
rect 11442 8878 11454 8930
rect 11506 8878 11518 8930
rect 13346 8878 13358 8930
rect 13410 8878 13422 8930
rect 16146 8878 16158 8930
rect 16210 8878 16222 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 21410 8878 21422 8930
rect 21474 8878 21486 8930
rect 25330 8878 25342 8930
rect 25394 8878 25406 8930
rect 38210 8878 38222 8930
rect 38274 8878 38286 8930
rect 41122 8878 41134 8930
rect 41186 8878 41198 8930
rect 7422 8866 7474 8878
rect 20526 8866 20578 8878
rect 34638 8866 34690 8878
rect 42814 8866 42866 8878
rect 44718 8930 44770 8942
rect 52546 8878 52558 8930
rect 52610 8878 52622 8930
rect 44718 8866 44770 8878
rect 10558 8818 10610 8830
rect 19518 8818 19570 8830
rect 16706 8766 16718 8818
rect 16770 8766 16782 8818
rect 18050 8766 18062 8818
rect 18114 8766 18126 8818
rect 10558 8754 10610 8766
rect 19518 8754 19570 8766
rect 22542 8818 22594 8830
rect 22542 8754 22594 8766
rect 43934 8818 43986 8830
rect 43934 8754 43986 8766
rect 44270 8818 44322 8830
rect 44270 8754 44322 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 19294 8482 19346 8494
rect 19294 8418 19346 8430
rect 19966 8482 20018 8494
rect 19966 8418 20018 8430
rect 44942 8482 44994 8494
rect 44942 8418 44994 8430
rect 9550 8370 9602 8382
rect 19070 8370 19122 8382
rect 37438 8370 37490 8382
rect 6290 8318 6302 8370
rect 6354 8318 6366 8370
rect 11890 8318 11902 8370
rect 11954 8318 11966 8370
rect 12786 8318 12798 8370
rect 12850 8318 12862 8370
rect 14690 8318 14702 8370
rect 14754 8318 14766 8370
rect 20626 8318 20638 8370
rect 20690 8318 20702 8370
rect 24882 8318 24894 8370
rect 24946 8318 24958 8370
rect 28466 8318 28478 8370
rect 28530 8318 28542 8370
rect 30930 8318 30942 8370
rect 30994 8318 31006 8370
rect 9550 8306 9602 8318
rect 19070 8306 19122 8318
rect 37438 8306 37490 8318
rect 37998 8370 38050 8382
rect 37998 8306 38050 8318
rect 41246 8370 41298 8382
rect 41246 8306 41298 8318
rect 45278 8370 45330 8382
rect 45278 8306 45330 8318
rect 57934 8370 57986 8382
rect 57934 8306 57986 8318
rect 6750 8258 6802 8270
rect 8430 8258 8482 8270
rect 11230 8258 11282 8270
rect 13358 8258 13410 8270
rect 7186 8206 7198 8258
rect 7250 8206 7262 8258
rect 8866 8206 8878 8258
rect 8930 8206 8942 8258
rect 12226 8206 12238 8258
rect 12290 8206 12302 8258
rect 13010 8206 13022 8258
rect 13074 8206 13086 8258
rect 6750 8194 6802 8206
rect 8430 8194 8482 8206
rect 11230 8194 11282 8206
rect 13358 8194 13410 8206
rect 13694 8258 13746 8270
rect 18734 8258 18786 8270
rect 14578 8206 14590 8258
rect 14642 8206 14654 8258
rect 14914 8206 14926 8258
rect 14978 8206 14990 8258
rect 16482 8206 16494 8258
rect 16546 8206 16558 8258
rect 17714 8206 17726 8258
rect 17778 8206 17790 8258
rect 13694 8194 13746 8206
rect 18734 8194 18786 8206
rect 19518 8258 19570 8270
rect 19518 8194 19570 8206
rect 21982 8258 22034 8270
rect 21982 8194 22034 8206
rect 22542 8258 22594 8270
rect 22542 8194 22594 8206
rect 23102 8258 23154 8270
rect 25790 8258 25842 8270
rect 29374 8258 29426 8270
rect 24210 8206 24222 8258
rect 24274 8206 24286 8258
rect 27682 8206 27694 8258
rect 27746 8206 27758 8258
rect 28018 8206 28030 8258
rect 28082 8206 28094 8258
rect 23102 8194 23154 8206
rect 25790 8194 25842 8206
rect 29374 8194 29426 8206
rect 29934 8258 29986 8270
rect 37102 8258 37154 8270
rect 32386 8206 32398 8258
rect 32450 8206 32462 8258
rect 33618 8206 33630 8258
rect 33682 8206 33694 8258
rect 35634 8206 35646 8258
rect 35698 8206 35710 8258
rect 29934 8194 29986 8206
rect 37102 8194 37154 8206
rect 40350 8258 40402 8270
rect 45054 8258 45106 8270
rect 40562 8206 40574 8258
rect 40626 8206 40638 8258
rect 40350 8194 40402 8206
rect 45054 8194 45106 8206
rect 47742 8258 47794 8270
rect 47742 8194 47794 8206
rect 47854 8258 47906 8270
rect 47854 8194 47906 8206
rect 47966 8258 48018 8270
rect 47966 8194 48018 8206
rect 48638 8258 48690 8270
rect 48638 8194 48690 8206
rect 48974 8258 49026 8270
rect 48974 8194 49026 8206
rect 49310 8258 49362 8270
rect 55570 8206 55582 8258
rect 55634 8206 55646 8258
rect 49310 8194 49362 8206
rect 7646 8146 7698 8158
rect 7646 8082 7698 8094
rect 13582 8146 13634 8158
rect 20190 8146 20242 8158
rect 14466 8094 14478 8146
rect 14530 8094 14542 8146
rect 16370 8094 16382 8146
rect 16434 8094 16446 8146
rect 13582 8082 13634 8094
rect 20190 8082 20242 8094
rect 21646 8146 21698 8158
rect 26350 8146 26402 8158
rect 30606 8146 30658 8158
rect 24546 8094 24558 8146
rect 24610 8094 24622 8146
rect 28130 8094 28142 8146
rect 28194 8094 28206 8146
rect 21646 8082 21698 8094
rect 26350 8082 26402 8094
rect 30606 8082 30658 8094
rect 30830 8146 30882 8158
rect 36318 8146 36370 8158
rect 31938 8094 31950 8146
rect 32002 8094 32014 8146
rect 34066 8094 34078 8146
rect 34130 8094 34142 8146
rect 30830 8082 30882 8094
rect 36318 8082 36370 8094
rect 37214 8146 37266 8158
rect 37214 8082 37266 8094
rect 37550 8146 37602 8158
rect 37550 8082 37602 8094
rect 38446 8146 38498 8158
rect 38446 8082 38498 8094
rect 45390 8146 45442 8158
rect 45390 8082 45442 8094
rect 45726 8146 45778 8158
rect 45726 8082 45778 8094
rect 45950 8146 46002 8158
rect 45950 8082 46002 8094
rect 46286 8146 46338 8158
rect 46286 8082 46338 8094
rect 8206 8034 8258 8046
rect 8206 7970 8258 7982
rect 9886 8034 9938 8046
rect 9886 7970 9938 7982
rect 10334 8034 10386 8046
rect 10334 7970 10386 7982
rect 10670 8034 10722 8046
rect 26798 8034 26850 8046
rect 30382 8034 30434 8046
rect 34974 8034 35026 8046
rect 46174 8034 46226 8046
rect 48862 8034 48914 8046
rect 17602 7982 17614 8034
rect 17666 7982 17678 8034
rect 27234 7982 27246 8034
rect 27298 7982 27310 8034
rect 33394 7982 33406 8034
rect 33458 7982 33470 8034
rect 35858 7982 35870 8034
rect 35922 7982 35934 8034
rect 48402 7982 48414 8034
rect 48466 7982 48478 8034
rect 10670 7970 10722 7982
rect 26798 7970 26850 7982
rect 30382 7970 30434 7982
rect 34974 7970 35026 7982
rect 46174 7970 46226 7982
rect 48862 7970 48914 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 6862 7698 6914 7710
rect 6862 7634 6914 7646
rect 7982 7698 8034 7710
rect 7982 7634 8034 7646
rect 9102 7698 9154 7710
rect 9102 7634 9154 7646
rect 15934 7698 15986 7710
rect 15934 7634 15986 7646
rect 17614 7698 17666 7710
rect 17614 7634 17666 7646
rect 17950 7698 18002 7710
rect 20302 7698 20354 7710
rect 19058 7646 19070 7698
rect 19122 7646 19134 7698
rect 17950 7634 18002 7646
rect 20302 7634 20354 7646
rect 35086 7698 35138 7710
rect 36642 7646 36654 7698
rect 36706 7646 36718 7698
rect 51538 7646 51550 7698
rect 51602 7646 51614 7698
rect 35086 7634 35138 7646
rect 13806 7586 13858 7598
rect 15710 7586 15762 7598
rect 12674 7534 12686 7586
rect 12738 7534 12750 7586
rect 15474 7534 15486 7586
rect 15538 7534 15550 7586
rect 13806 7522 13858 7534
rect 15710 7522 15762 7534
rect 16830 7586 16882 7598
rect 16830 7522 16882 7534
rect 17838 7586 17890 7598
rect 17838 7522 17890 7534
rect 20526 7586 20578 7598
rect 20526 7522 20578 7534
rect 20638 7586 20690 7598
rect 24670 7586 24722 7598
rect 23538 7534 23550 7586
rect 23602 7534 23614 7586
rect 20638 7522 20690 7534
rect 24670 7522 24722 7534
rect 25230 7586 25282 7598
rect 25230 7522 25282 7534
rect 25342 7586 25394 7598
rect 25342 7522 25394 7534
rect 26350 7586 26402 7598
rect 26350 7522 26402 7534
rect 35534 7586 35586 7598
rect 35534 7522 35586 7534
rect 38446 7586 38498 7598
rect 50642 7534 50654 7586
rect 50706 7534 50718 7586
rect 38446 7522 38498 7534
rect 9550 7474 9602 7486
rect 9550 7410 9602 7422
rect 10110 7474 10162 7486
rect 13358 7474 13410 7486
rect 11778 7422 11790 7474
rect 11842 7422 11854 7474
rect 10110 7410 10162 7422
rect 13358 7410 13410 7422
rect 13470 7474 13522 7486
rect 16046 7474 16098 7486
rect 14130 7422 14142 7474
rect 14194 7422 14206 7474
rect 15138 7422 15150 7474
rect 15202 7422 15214 7474
rect 13470 7410 13522 7422
rect 16046 7410 16098 7422
rect 17278 7474 17330 7486
rect 17278 7410 17330 7422
rect 22094 7474 22146 7486
rect 22094 7410 22146 7422
rect 22654 7474 22706 7486
rect 32286 7474 32338 7486
rect 23202 7422 23214 7474
rect 23266 7422 23278 7474
rect 24434 7422 24446 7474
rect 24498 7422 24510 7474
rect 25890 7422 25902 7474
rect 25954 7422 25966 7474
rect 27234 7422 27246 7474
rect 27298 7422 27310 7474
rect 29138 7422 29150 7474
rect 29202 7422 29214 7474
rect 30370 7422 30382 7474
rect 30434 7422 30446 7474
rect 30818 7422 30830 7474
rect 30882 7422 30894 7474
rect 31714 7422 31726 7474
rect 31778 7422 31790 7474
rect 22654 7410 22706 7422
rect 32286 7410 32338 7422
rect 33182 7474 33234 7486
rect 33182 7410 33234 7422
rect 33742 7474 33794 7486
rect 33742 7410 33794 7422
rect 34078 7474 34130 7486
rect 34078 7410 34130 7422
rect 34302 7474 34354 7486
rect 34302 7410 34354 7422
rect 34750 7474 34802 7486
rect 37886 7474 37938 7486
rect 44606 7474 44658 7486
rect 48862 7474 48914 7486
rect 37314 7422 37326 7474
rect 37378 7422 37390 7474
rect 38658 7422 38670 7474
rect 38722 7422 38734 7474
rect 39330 7422 39342 7474
rect 39394 7422 39406 7474
rect 41122 7422 41134 7474
rect 41186 7422 41198 7474
rect 43922 7422 43934 7474
rect 43986 7422 43998 7474
rect 45490 7422 45502 7474
rect 45554 7422 45566 7474
rect 34750 7410 34802 7422
rect 37886 7410 37938 7422
rect 44606 7410 44658 7422
rect 48862 7410 48914 7422
rect 48974 7474 49026 7486
rect 48974 7410 49026 7422
rect 49310 7474 49362 7486
rect 50530 7422 50542 7474
rect 50594 7422 50606 7474
rect 51426 7422 51438 7474
rect 51490 7422 51502 7474
rect 49310 7410 49362 7422
rect 7198 7362 7250 7374
rect 7198 7298 7250 7310
rect 7758 7362 7810 7374
rect 7758 7298 7810 7310
rect 8542 7362 8594 7374
rect 8542 7298 8594 7310
rect 10782 7362 10834 7374
rect 18510 7362 18562 7374
rect 11330 7310 11342 7362
rect 11394 7310 11406 7362
rect 14690 7310 14702 7362
rect 14754 7310 14766 7362
rect 10782 7298 10834 7310
rect 18510 7298 18562 7310
rect 19742 7362 19794 7374
rect 19742 7298 19794 7310
rect 21310 7362 21362 7374
rect 21310 7298 21362 7310
rect 21758 7362 21810 7374
rect 34190 7362 34242 7374
rect 23426 7310 23438 7362
rect 23490 7310 23502 7362
rect 27794 7310 27806 7362
rect 27858 7310 27870 7362
rect 29026 7310 29038 7362
rect 29090 7310 29102 7362
rect 30706 7310 30718 7362
rect 30770 7310 30782 7362
rect 21758 7298 21810 7310
rect 34190 7298 34242 7310
rect 35646 7362 35698 7374
rect 35646 7298 35698 7310
rect 36094 7362 36146 7374
rect 36094 7298 36146 7310
rect 37998 7362 38050 7374
rect 37998 7298 38050 7310
rect 39566 7362 39618 7374
rect 39566 7298 39618 7310
rect 39678 7362 39730 7374
rect 39678 7298 39730 7310
rect 40126 7362 40178 7374
rect 41570 7310 41582 7362
rect 41634 7310 41646 7362
rect 46050 7310 46062 7362
rect 46114 7310 46126 7362
rect 40126 7298 40178 7310
rect 13694 7250 13746 7262
rect 7186 7198 7198 7250
rect 7250 7247 7262 7250
rect 7410 7247 7422 7250
rect 7250 7201 7422 7247
rect 7250 7198 7262 7201
rect 7410 7198 7422 7201
rect 7474 7198 7486 7250
rect 13694 7186 13746 7198
rect 18734 7250 18786 7262
rect 18734 7186 18786 7198
rect 20638 7250 20690 7262
rect 20638 7186 20690 7198
rect 25342 7250 25394 7262
rect 35758 7250 35810 7262
rect 31938 7198 31950 7250
rect 32002 7198 32014 7250
rect 25342 7186 25394 7198
rect 35758 7186 35810 7198
rect 36318 7250 36370 7262
rect 36318 7186 36370 7198
rect 38334 7250 38386 7262
rect 49198 7250 49250 7262
rect 41906 7198 41918 7250
rect 41970 7198 41982 7250
rect 38334 7186 38386 7198
rect 49198 7186 49250 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 8206 6914 8258 6926
rect 15598 6914 15650 6926
rect 6850 6862 6862 6914
rect 6914 6911 6926 6914
rect 7298 6911 7310 6914
rect 6914 6865 7310 6911
rect 6914 6862 6926 6865
rect 7298 6862 7310 6865
rect 7362 6862 7374 6914
rect 14018 6862 14030 6914
rect 14082 6862 14094 6914
rect 35522 6862 35534 6914
rect 35586 6911 35598 6914
rect 36530 6911 36542 6914
rect 35586 6865 36542 6911
rect 35586 6862 35598 6865
rect 36530 6862 36542 6865
rect 36594 6862 36606 6914
rect 45826 6862 45838 6914
rect 45890 6862 45902 6914
rect 8206 6850 8258 6862
rect 15598 6850 15650 6862
rect 7310 6802 7362 6814
rect 7310 6738 7362 6750
rect 7646 6802 7698 6814
rect 7646 6738 7698 6750
rect 7982 6802 8034 6814
rect 22542 6802 22594 6814
rect 15922 6750 15934 6802
rect 15986 6750 15998 6802
rect 20178 6750 20190 6802
rect 20242 6750 20254 6802
rect 7982 6738 8034 6750
rect 22542 6738 22594 6750
rect 27806 6802 27858 6814
rect 36206 6802 36258 6814
rect 29474 6750 29486 6802
rect 29538 6750 29550 6802
rect 37090 6750 37102 6802
rect 37154 6750 37166 6802
rect 40786 6750 40798 6802
rect 40850 6750 40862 6802
rect 45154 6750 45166 6802
rect 45218 6750 45230 6802
rect 47730 6750 47742 6802
rect 47794 6750 47806 6802
rect 50530 6750 50542 6802
rect 50594 6750 50606 6802
rect 27806 6738 27858 6750
rect 36206 6738 36258 6750
rect 9326 6690 9378 6702
rect 9326 6626 9378 6638
rect 10222 6690 10274 6702
rect 10222 6626 10274 6638
rect 10782 6690 10834 6702
rect 10782 6626 10834 6638
rect 11118 6690 11170 6702
rect 12910 6690 12962 6702
rect 16158 6690 16210 6702
rect 11778 6638 11790 6690
rect 11842 6638 11854 6690
rect 13570 6638 13582 6690
rect 13634 6638 13646 6690
rect 14018 6638 14030 6690
rect 14082 6638 14094 6690
rect 14914 6638 14926 6690
rect 14978 6638 14990 6690
rect 11118 6626 11170 6638
rect 12910 6626 12962 6638
rect 16158 6626 16210 6638
rect 16606 6690 16658 6702
rect 18398 6690 18450 6702
rect 17490 6638 17502 6690
rect 17554 6638 17566 6690
rect 16606 6626 16658 6638
rect 18398 6626 18450 6638
rect 18958 6690 19010 6702
rect 28254 6690 28306 6702
rect 29934 6690 29986 6702
rect 35198 6690 35250 6702
rect 37998 6690 38050 6702
rect 42814 6690 42866 6702
rect 19282 6638 19294 6690
rect 19346 6638 19358 6690
rect 19842 6638 19854 6690
rect 19906 6638 19918 6690
rect 21410 6638 21422 6690
rect 21474 6638 21486 6690
rect 22978 6638 22990 6690
rect 23042 6638 23054 6690
rect 24658 6638 24670 6690
rect 24722 6638 24734 6690
rect 26226 6638 26238 6690
rect 26290 6638 26302 6690
rect 29362 6638 29374 6690
rect 29426 6638 29438 6690
rect 30818 6638 30830 6690
rect 30882 6638 30894 6690
rect 32274 6638 32286 6690
rect 32338 6638 32350 6690
rect 34066 6638 34078 6690
rect 34130 6638 34142 6690
rect 37314 6638 37326 6690
rect 37378 6638 37390 6690
rect 40898 6638 40910 6690
rect 40962 6638 40974 6690
rect 41346 6638 41358 6690
rect 41410 6638 41422 6690
rect 42578 6638 42590 6690
rect 42642 6638 42654 6690
rect 18958 6626 19010 6638
rect 28254 6626 28306 6638
rect 29934 6626 29986 6638
rect 35198 6626 35250 6638
rect 37998 6626 38050 6638
rect 42814 6626 42866 6638
rect 43486 6690 43538 6702
rect 49870 6690 49922 6702
rect 45266 6638 45278 6690
rect 45330 6638 45342 6690
rect 49410 6638 49422 6690
rect 49474 6638 49486 6690
rect 50642 6638 50654 6690
rect 50706 6638 50718 6690
rect 43486 6626 43538 6638
rect 49870 6626 49922 6638
rect 9886 6578 9938 6590
rect 9886 6514 9938 6526
rect 16830 6578 16882 6590
rect 28590 6578 28642 6590
rect 38446 6578 38498 6590
rect 20066 6526 20078 6578
rect 20130 6526 20142 6578
rect 21522 6526 21534 6578
rect 21586 6526 21598 6578
rect 22082 6526 22094 6578
rect 22146 6526 22158 6578
rect 22754 6526 22766 6578
rect 22818 6526 22830 6578
rect 26114 6526 26126 6578
rect 26178 6526 26190 6578
rect 30594 6526 30606 6578
rect 30658 6526 30670 6578
rect 34738 6526 34750 6578
rect 34802 6526 34814 6578
rect 16830 6514 16882 6526
rect 28590 6514 28642 6526
rect 38446 6514 38498 6526
rect 41918 6578 41970 6590
rect 51326 6578 51378 6590
rect 47954 6526 47966 6578
rect 48018 6526 48030 6578
rect 41918 6514 41970 6526
rect 51326 6514 51378 6526
rect 51662 6578 51714 6590
rect 51662 6514 51714 6526
rect 8990 6466 9042 6478
rect 8530 6414 8542 6466
rect 8594 6414 8606 6466
rect 8990 6402 9042 6414
rect 15262 6466 15314 6478
rect 15262 6402 15314 6414
rect 15822 6466 15874 6478
rect 15822 6402 15874 6414
rect 16494 6466 16546 6478
rect 27246 6466 27298 6478
rect 26674 6414 26686 6466
rect 26738 6414 26750 6466
rect 16494 6402 16546 6414
rect 27246 6402 27298 6414
rect 28478 6466 28530 6478
rect 35646 6466 35698 6478
rect 34514 6414 34526 6466
rect 34578 6414 34590 6466
rect 28478 6402 28530 6414
rect 35646 6402 35698 6414
rect 39118 6466 39170 6478
rect 51986 6414 51998 6466
rect 52050 6414 52062 6466
rect 39118 6402 39170 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 7758 6130 7810 6142
rect 7758 6066 7810 6078
rect 8094 6130 8146 6142
rect 8094 6066 8146 6078
rect 8430 6130 8482 6142
rect 8430 6066 8482 6078
rect 9774 6130 9826 6142
rect 9774 6066 9826 6078
rect 11230 6130 11282 6142
rect 11230 6066 11282 6078
rect 11678 6130 11730 6142
rect 11678 6066 11730 6078
rect 12238 6130 12290 6142
rect 16046 6130 16098 6142
rect 12786 6078 12798 6130
rect 12850 6078 12862 6130
rect 12238 6066 12290 6078
rect 16046 6066 16098 6078
rect 19406 6130 19458 6142
rect 27806 6130 27858 6142
rect 26786 6078 26798 6130
rect 26850 6078 26862 6130
rect 19406 6066 19458 6078
rect 27806 6066 27858 6078
rect 35982 6130 36034 6142
rect 35982 6066 36034 6078
rect 36542 6130 36594 6142
rect 36542 6066 36594 6078
rect 37326 6130 37378 6142
rect 37326 6066 37378 6078
rect 46734 6130 46786 6142
rect 46734 6066 46786 6078
rect 47294 6130 47346 6142
rect 47294 6066 47346 6078
rect 10670 6018 10722 6030
rect 10670 5954 10722 5966
rect 14478 6018 14530 6030
rect 14478 5954 14530 5966
rect 15262 6018 15314 6030
rect 15262 5954 15314 5966
rect 18062 6018 18114 6030
rect 18062 5954 18114 5966
rect 19182 6018 19234 6030
rect 19182 5954 19234 5966
rect 24558 6018 24610 6030
rect 27358 6018 27410 6030
rect 32174 6018 32226 6030
rect 40238 6018 40290 6030
rect 25218 5966 25230 6018
rect 25282 5966 25294 6018
rect 27570 5966 27582 6018
rect 27634 5966 27646 6018
rect 30146 5966 30158 6018
rect 30210 5966 30222 6018
rect 30594 5966 30606 6018
rect 30658 5966 30670 6018
rect 33618 5966 33630 6018
rect 33682 5966 33694 6018
rect 35186 5966 35198 6018
rect 35250 5966 35262 6018
rect 24558 5954 24610 5966
rect 27358 5954 27410 5966
rect 32174 5954 32226 5966
rect 40238 5954 40290 5966
rect 46510 6018 46562 6030
rect 46510 5954 46562 5966
rect 47182 6018 47234 6030
rect 47182 5954 47234 5966
rect 13694 5906 13746 5918
rect 10210 5854 10222 5906
rect 10274 5854 10286 5906
rect 12562 5854 12574 5906
rect 12626 5854 12638 5906
rect 13234 5854 13246 5906
rect 13298 5854 13310 5906
rect 13694 5842 13746 5854
rect 13918 5906 13970 5918
rect 14702 5906 14754 5918
rect 17390 5906 17442 5918
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 15026 5854 15038 5906
rect 15090 5854 15102 5906
rect 13918 5842 13970 5854
rect 14702 5842 14754 5854
rect 17390 5842 17442 5854
rect 17838 5906 17890 5918
rect 17838 5842 17890 5854
rect 19070 5906 19122 5918
rect 28142 5906 28194 5918
rect 31950 5906 32002 5918
rect 20178 5854 20190 5906
rect 20242 5854 20254 5906
rect 21298 5854 21310 5906
rect 21362 5854 21374 5906
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 23090 5854 23102 5906
rect 23154 5854 23166 5906
rect 26226 5854 26238 5906
rect 26290 5854 26302 5906
rect 28802 5854 28814 5906
rect 28866 5854 28878 5906
rect 29922 5854 29934 5906
rect 29986 5854 29998 5906
rect 31154 5854 31166 5906
rect 31218 5854 31230 5906
rect 31490 5854 31502 5906
rect 31554 5854 31566 5906
rect 19070 5842 19122 5854
rect 28142 5842 28194 5854
rect 31950 5842 32002 5854
rect 32286 5906 32338 5918
rect 40126 5906 40178 5918
rect 42366 5906 42418 5918
rect 34066 5854 34078 5906
rect 34130 5854 34142 5906
rect 34962 5854 34974 5906
rect 35026 5854 35038 5906
rect 39778 5854 39790 5906
rect 39842 5854 39854 5906
rect 42018 5854 42030 5906
rect 42082 5854 42094 5906
rect 32286 5842 32338 5854
rect 40126 5842 40178 5854
rect 42366 5842 42418 5854
rect 42590 5906 42642 5918
rect 42590 5842 42642 5854
rect 47518 5906 47570 5918
rect 47518 5842 47570 5854
rect 8990 5794 9042 5806
rect 8990 5730 9042 5742
rect 14142 5794 14194 5806
rect 14142 5730 14194 5742
rect 16382 5794 16434 5806
rect 16382 5730 16434 5742
rect 16830 5794 16882 5806
rect 16830 5730 16882 5742
rect 17614 5794 17666 5806
rect 17614 5730 17666 5742
rect 18846 5794 18898 5806
rect 18846 5730 18898 5742
rect 19742 5794 19794 5806
rect 30046 5794 30098 5806
rect 36878 5794 36930 5806
rect 27234 5742 27246 5794
rect 27298 5742 27310 5794
rect 30818 5742 30830 5794
rect 30882 5742 30894 5794
rect 19742 5730 19794 5742
rect 30046 5730 30098 5742
rect 36878 5730 36930 5742
rect 46622 5794 46674 5806
rect 46622 5730 46674 5742
rect 15374 5682 15426 5694
rect 28254 5682 28306 5694
rect 15922 5630 15934 5682
rect 15986 5679 15998 5682
rect 16370 5679 16382 5682
rect 15986 5633 16382 5679
rect 15986 5630 15998 5633
rect 16370 5630 16382 5633
rect 16434 5630 16446 5682
rect 23426 5630 23438 5682
rect 23490 5630 23502 5682
rect 15374 5618 15426 5630
rect 28254 5618 28306 5630
rect 39454 5682 39506 5694
rect 39454 5618 39506 5630
rect 39790 5682 39842 5694
rect 39790 5618 39842 5630
rect 58158 5682 58210 5694
rect 58158 5618 58210 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 13470 5346 13522 5358
rect 13470 5282 13522 5294
rect 16942 5346 16994 5358
rect 16942 5282 16994 5294
rect 21422 5346 21474 5358
rect 27682 5294 27694 5346
rect 27746 5294 27758 5346
rect 31602 5294 31614 5346
rect 31666 5294 31678 5346
rect 21422 5282 21474 5294
rect 9214 5234 9266 5246
rect 9214 5170 9266 5182
rect 9662 5234 9714 5246
rect 9662 5170 9714 5182
rect 10110 5234 10162 5246
rect 13694 5234 13746 5246
rect 11554 5182 11566 5234
rect 11618 5182 11630 5234
rect 10110 5170 10162 5182
rect 13694 5170 13746 5182
rect 15150 5234 15202 5246
rect 15150 5170 15202 5182
rect 16718 5234 16770 5246
rect 26574 5234 26626 5246
rect 22530 5182 22542 5234
rect 22594 5182 22606 5234
rect 24882 5182 24894 5234
rect 24946 5182 24958 5234
rect 16718 5170 16770 5182
rect 26574 5170 26626 5182
rect 27134 5234 27186 5246
rect 27134 5170 27186 5182
rect 27358 5234 27410 5246
rect 32062 5234 32114 5246
rect 28466 5182 28478 5234
rect 28530 5182 28542 5234
rect 27358 5170 27410 5182
rect 32062 5170 32114 5182
rect 33294 5234 33346 5246
rect 33294 5170 33346 5182
rect 34302 5234 34354 5246
rect 34302 5170 34354 5182
rect 35086 5234 35138 5246
rect 35086 5170 35138 5182
rect 35422 5234 35474 5246
rect 58158 5234 58210 5246
rect 38882 5182 38894 5234
rect 38946 5182 38958 5234
rect 41122 5182 41134 5234
rect 41186 5182 41198 5234
rect 45490 5182 45502 5234
rect 45554 5182 45566 5234
rect 35422 5170 35474 5182
rect 58158 5170 58210 5182
rect 10334 5122 10386 5134
rect 10334 5058 10386 5070
rect 11118 5122 11170 5134
rect 11118 5058 11170 5070
rect 12238 5122 12290 5134
rect 12238 5058 12290 5070
rect 14030 5122 14082 5134
rect 14030 5058 14082 5070
rect 14926 5122 14978 5134
rect 14926 5058 14978 5070
rect 15374 5122 15426 5134
rect 15374 5058 15426 5070
rect 15598 5122 15650 5134
rect 15598 5058 15650 5070
rect 16270 5122 16322 5134
rect 16270 5058 16322 5070
rect 16606 5122 16658 5134
rect 16606 5058 16658 5070
rect 18286 5122 18338 5134
rect 18286 5058 18338 5070
rect 19070 5122 19122 5134
rect 20862 5122 20914 5134
rect 32398 5122 32450 5134
rect 20290 5070 20302 5122
rect 20354 5070 20366 5122
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 22754 5070 22766 5122
rect 22818 5070 22830 5122
rect 24434 5070 24446 5122
rect 24498 5070 24510 5122
rect 26002 5070 26014 5122
rect 26066 5070 26078 5122
rect 28130 5070 28142 5122
rect 28194 5070 28206 5122
rect 29138 5070 29150 5122
rect 29202 5070 29214 5122
rect 30818 5070 30830 5122
rect 30882 5070 30894 5122
rect 32162 5070 32174 5122
rect 32226 5070 32238 5122
rect 19070 5058 19122 5070
rect 20862 5058 20914 5070
rect 32398 5058 32450 5070
rect 33742 5122 33794 5134
rect 39790 5122 39842 5134
rect 43374 5122 43426 5134
rect 39330 5070 39342 5122
rect 39394 5070 39406 5122
rect 40114 5070 40126 5122
rect 40178 5070 40190 5122
rect 40674 5070 40686 5122
rect 40738 5070 40750 5122
rect 42802 5070 42814 5122
rect 42866 5070 42878 5122
rect 33742 5058 33794 5070
rect 39790 5058 39842 5070
rect 43374 5058 43426 5070
rect 43486 5122 43538 5134
rect 43486 5058 43538 5070
rect 43822 5122 43874 5134
rect 43822 5058 43874 5070
rect 45166 5122 45218 5134
rect 48078 5122 48130 5134
rect 46722 5070 46734 5122
rect 46786 5070 46798 5122
rect 47394 5070 47406 5122
rect 47458 5070 47470 5122
rect 48626 5070 48638 5122
rect 48690 5070 48702 5122
rect 45166 5058 45218 5070
rect 48078 5058 48130 5070
rect 18510 5010 18562 5022
rect 26350 5010 26402 5022
rect 45390 5010 45442 5022
rect 10658 4958 10670 5010
rect 10722 4958 10734 5010
rect 17490 4958 17502 5010
rect 17554 4958 17566 5010
rect 21410 4958 21422 5010
rect 21474 4958 21486 5010
rect 30034 4958 30046 5010
rect 30098 4958 30110 5010
rect 41234 4958 41246 5010
rect 41298 4958 41310 5010
rect 46162 4958 46174 5010
rect 46226 4958 46238 5010
rect 18510 4946 18562 4958
rect 26350 4946 26402 4958
rect 45390 4946 45442 4958
rect 13918 4898 13970 4910
rect 12562 4846 12574 4898
rect 12626 4846 12638 4898
rect 13918 4834 13970 4846
rect 14142 4898 14194 4910
rect 14142 4834 14194 4846
rect 14814 4898 14866 4910
rect 14814 4834 14866 4846
rect 18062 4898 18114 4910
rect 18062 4834 18114 4846
rect 18174 4898 18226 4910
rect 18174 4834 18226 4846
rect 26462 4898 26514 4910
rect 26462 4834 26514 4846
rect 26686 4898 26738 4910
rect 26686 4834 26738 4846
rect 44158 4898 44210 4910
rect 44158 4834 44210 4846
rect 48414 4898 48466 4910
rect 48414 4834 48466 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 10670 4562 10722 4574
rect 10670 4498 10722 4510
rect 11230 4562 11282 4574
rect 11230 4498 11282 4510
rect 13694 4562 13746 4574
rect 13694 4498 13746 4510
rect 16046 4562 16098 4574
rect 16046 4498 16098 4510
rect 17726 4562 17778 4574
rect 17726 4498 17778 4510
rect 24782 4562 24834 4574
rect 24782 4498 24834 4510
rect 27246 4562 27298 4574
rect 27246 4498 27298 4510
rect 28366 4562 28418 4574
rect 28366 4498 28418 4510
rect 29150 4562 29202 4574
rect 33182 4562 33234 4574
rect 31602 4510 31614 4562
rect 31666 4510 31678 4562
rect 29150 4498 29202 4510
rect 33182 4498 33234 4510
rect 34190 4562 34242 4574
rect 34190 4498 34242 4510
rect 34526 4562 34578 4574
rect 34526 4498 34578 4510
rect 11902 4450 11954 4462
rect 11902 4386 11954 4398
rect 12238 4450 12290 4462
rect 12238 4386 12290 4398
rect 17614 4450 17666 4462
rect 17614 4386 17666 4398
rect 17950 4450 18002 4462
rect 17950 4386 18002 4398
rect 18846 4450 18898 4462
rect 18846 4386 18898 4398
rect 25230 4450 25282 4462
rect 40910 4450 40962 4462
rect 58158 4450 58210 4462
rect 30930 4398 30942 4450
rect 30994 4398 31006 4450
rect 46274 4398 46286 4450
rect 46338 4398 46350 4450
rect 25230 4386 25282 4398
rect 40910 4386 40962 4398
rect 58158 4386 58210 4398
rect 13358 4338 13410 4350
rect 12898 4286 12910 4338
rect 12962 4286 12974 4338
rect 13358 4274 13410 4286
rect 14254 4338 14306 4350
rect 16270 4338 16322 4350
rect 14802 4286 14814 4338
rect 14866 4286 14878 4338
rect 14254 4274 14306 4286
rect 16270 4274 16322 4286
rect 18062 4338 18114 4350
rect 18062 4274 18114 4286
rect 19294 4338 19346 4350
rect 21534 4338 21586 4350
rect 25790 4338 25842 4350
rect 27806 4338 27858 4350
rect 19954 4286 19966 4338
rect 20018 4286 20030 4338
rect 21746 4286 21758 4338
rect 21810 4286 21822 4338
rect 23426 4286 23438 4338
rect 23490 4286 23502 4338
rect 26450 4286 26462 4338
rect 26514 4286 26526 4338
rect 19294 4274 19346 4286
rect 21534 4274 21586 4286
rect 25790 4274 25842 4286
rect 27806 4274 27858 4286
rect 28590 4338 28642 4350
rect 28590 4274 28642 4286
rect 29486 4338 29538 4350
rect 40350 4338 40402 4350
rect 47742 4338 47794 4350
rect 30594 4286 30606 4338
rect 30658 4286 30670 4338
rect 31490 4286 31502 4338
rect 31554 4286 31566 4338
rect 39666 4286 39678 4338
rect 39730 4286 39742 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 29486 4274 29538 4286
rect 40350 4274 40402 4286
rect 47742 4274 47794 4286
rect 10334 4226 10386 4238
rect 10334 4162 10386 4174
rect 11678 4226 11730 4238
rect 11678 4162 11730 4174
rect 15262 4226 15314 4238
rect 18958 4226 19010 4238
rect 32174 4226 32226 4238
rect 16706 4174 16718 4226
rect 16770 4174 16782 4226
rect 20962 4174 20974 4226
rect 21026 4174 21038 4226
rect 26786 4174 26798 4226
rect 26850 4174 26862 4226
rect 29922 4174 29934 4226
rect 29986 4174 29998 4226
rect 15262 4162 15314 4174
rect 18958 4162 19010 4174
rect 32174 4162 32226 4174
rect 33630 4226 33682 4238
rect 39890 4174 39902 4226
rect 39954 4174 39966 4226
rect 46498 4174 46510 4226
rect 46562 4174 46574 4226
rect 33630 4162 33682 4174
rect 19182 4114 19234 4126
rect 47854 4114 47906 4126
rect 22978 4062 22990 4114
rect 23042 4062 23054 4114
rect 46610 4062 46622 4114
rect 46674 4062 46686 4114
rect 19182 4050 19234 4062
rect 47854 4050 47906 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 25790 3778 25842 3790
rect 10322 3726 10334 3778
rect 10386 3775 10398 3778
rect 12674 3775 12686 3778
rect 10386 3729 12686 3775
rect 10386 3726 10398 3729
rect 12674 3726 12686 3729
rect 12738 3726 12750 3778
rect 25790 3714 25842 3726
rect 26126 3778 26178 3790
rect 28578 3726 28590 3778
rect 28642 3775 28654 3778
rect 29474 3775 29486 3778
rect 28642 3729 29486 3775
rect 28642 3726 28654 3729
rect 29474 3726 29486 3729
rect 29538 3726 29550 3778
rect 26126 3714 26178 3726
rect 6974 3666 7026 3678
rect 6974 3602 7026 3614
rect 10446 3666 10498 3678
rect 10446 3602 10498 3614
rect 10894 3666 10946 3678
rect 10894 3602 10946 3614
rect 11790 3666 11842 3678
rect 11790 3602 11842 3614
rect 12238 3666 12290 3678
rect 12238 3602 12290 3614
rect 12686 3666 12738 3678
rect 12686 3602 12738 3614
rect 13358 3666 13410 3678
rect 13358 3602 13410 3614
rect 13806 3666 13858 3678
rect 13806 3602 13858 3614
rect 14142 3666 14194 3678
rect 14142 3602 14194 3614
rect 16046 3666 16098 3678
rect 16046 3602 16098 3614
rect 16494 3666 16546 3678
rect 16494 3602 16546 3614
rect 17726 3666 17778 3678
rect 17726 3602 17778 3614
rect 18510 3666 18562 3678
rect 18510 3602 18562 3614
rect 18958 3666 19010 3678
rect 18958 3602 19010 3614
rect 19406 3666 19458 3678
rect 19406 3602 19458 3614
rect 20302 3666 20354 3678
rect 20302 3602 20354 3614
rect 21310 3666 21362 3678
rect 21310 3602 21362 3614
rect 21758 3666 21810 3678
rect 23998 3666 24050 3678
rect 22082 3614 22094 3666
rect 22146 3614 22158 3666
rect 21758 3602 21810 3614
rect 23998 3602 24050 3614
rect 25118 3666 25170 3678
rect 25118 3602 25170 3614
rect 27358 3666 27410 3678
rect 27358 3602 27410 3614
rect 28590 3666 28642 3678
rect 28590 3602 28642 3614
rect 29038 3666 29090 3678
rect 30830 3666 30882 3678
rect 30146 3614 30158 3666
rect 30210 3614 30222 3666
rect 29038 3602 29090 3614
rect 30830 3602 30882 3614
rect 31278 3666 31330 3678
rect 31278 3602 31330 3614
rect 33182 3666 33234 3678
rect 33182 3602 33234 3614
rect 33630 3666 33682 3678
rect 33630 3602 33682 3614
rect 34078 3666 34130 3678
rect 34078 3602 34130 3614
rect 49086 3666 49138 3678
rect 49086 3602 49138 3614
rect 52894 3666 52946 3678
rect 52894 3602 52946 3614
rect 15598 3554 15650 3566
rect 15598 3490 15650 3502
rect 17166 3554 17218 3566
rect 24558 3554 24610 3566
rect 27806 3554 27858 3566
rect 22418 3502 22430 3554
rect 22482 3502 22494 3554
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 26114 3502 26126 3554
rect 26178 3502 26190 3554
rect 26674 3502 26686 3554
rect 26738 3502 26750 3554
rect 17166 3490 17218 3502
rect 24558 3490 24610 3502
rect 27806 3490 27858 3502
rect 29710 3554 29762 3566
rect 29710 3490 29762 3502
rect 31614 3554 31666 3566
rect 40898 3502 40910 3554
rect 40962 3502 40974 3554
rect 44146 3502 44158 3554
rect 44210 3502 44222 3554
rect 48402 3502 48414 3554
rect 48466 3502 48478 3554
rect 52098 3502 52110 3554
rect 52162 3502 52174 3554
rect 31614 3490 31666 3502
rect 14590 3442 14642 3454
rect 14590 3378 14642 3390
rect 15150 3442 15202 3454
rect 15150 3378 15202 3390
rect 19854 3442 19906 3454
rect 19854 3378 19906 3390
rect 23214 3442 23266 3454
rect 23214 3378 23266 3390
rect 26462 3442 26514 3454
rect 26462 3378 26514 3390
rect 29486 3442 29538 3454
rect 29486 3378 29538 3390
rect 32398 3442 32450 3454
rect 32398 3378 32450 3390
rect 4846 3330 4898 3342
rect 4846 3266 4898 3278
rect 5630 3330 5682 3342
rect 5630 3266 5682 3278
rect 7646 3330 7698 3342
rect 7646 3266 7698 3278
rect 11342 3330 11394 3342
rect 11342 3266 11394 3278
rect 32734 3330 32786 3342
rect 32734 3266 32786 3278
rect 41470 3330 41522 3342
rect 41470 3266 41522 3278
rect 44942 3330 44994 3342
rect 44942 3266 44994 3278
rect 57710 3330 57762 3342
rect 57710 3266 57762 3278
rect 58158 3330 58210 3342
rect 58158 3266 58210 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 53790 56590 53842 56642
rect 55022 56590 55074 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 10334 56254 10386 56306
rect 11006 56254 11058 56306
rect 13694 56254 13746 56306
rect 25230 56254 25282 56306
rect 34302 56254 34354 56306
rect 48974 56254 49026 56306
rect 52222 56254 52274 56306
rect 54126 56254 54178 56306
rect 55022 56254 55074 56306
rect 55470 56254 55522 56306
rect 33742 56142 33794 56194
rect 25118 56030 25170 56082
rect 31166 56030 31218 56082
rect 32286 56030 32338 56082
rect 33294 56030 33346 56082
rect 33854 56030 33906 56082
rect 48190 56030 48242 56082
rect 51214 56030 51266 56082
rect 8318 55918 8370 55970
rect 19182 55918 19234 55970
rect 25790 55918 25842 55970
rect 26910 55918 26962 55970
rect 29598 55918 29650 55970
rect 33518 55918 33570 55970
rect 34750 55918 34802 55970
rect 55918 55918 55970 55970
rect 25230 55806 25282 55858
rect 58158 55806 58210 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 48190 55470 48242 55522
rect 29374 55358 29426 55410
rect 49646 55358 49698 55410
rect 53678 55358 53730 55410
rect 23774 55246 23826 55298
rect 29710 55246 29762 55298
rect 33070 55246 33122 55298
rect 33742 55246 33794 55298
rect 34078 55246 34130 55298
rect 35086 55246 35138 55298
rect 35422 55246 35474 55298
rect 36990 55246 37042 55298
rect 37214 55246 37266 55298
rect 39006 55246 39058 55298
rect 39566 55246 39618 55298
rect 40238 55246 40290 55298
rect 48750 55246 48802 55298
rect 51774 55246 51826 55298
rect 53006 55246 53058 55298
rect 19630 55134 19682 55186
rect 19966 55134 20018 55186
rect 20190 55134 20242 55186
rect 24894 55134 24946 55186
rect 25678 55134 25730 55186
rect 26462 55134 26514 55186
rect 27806 55134 27858 55186
rect 30830 55134 30882 55186
rect 32958 55134 33010 55186
rect 34526 55134 34578 55186
rect 37774 55134 37826 55186
rect 41022 55134 41074 55186
rect 42478 55134 42530 55186
rect 44830 55134 44882 55186
rect 45390 55134 45442 55186
rect 45502 55134 45554 55186
rect 45726 55134 45778 55186
rect 46846 55134 46898 55186
rect 46958 55134 47010 55186
rect 47070 55134 47122 55186
rect 47518 55134 47570 55186
rect 47854 55134 47906 55186
rect 57710 55134 57762 55186
rect 18734 55022 18786 55074
rect 19182 55022 19234 55074
rect 19854 55022 19906 55074
rect 20862 55022 20914 55074
rect 21310 55022 21362 55074
rect 21646 55022 21698 55074
rect 22206 55022 22258 55074
rect 22430 55022 22482 55074
rect 22766 55022 22818 55074
rect 25790 55022 25842 55074
rect 26014 55022 26066 55074
rect 26574 55022 26626 55074
rect 26798 55022 26850 55074
rect 27470 55022 27522 55074
rect 27918 55022 27970 55074
rect 28030 55022 28082 55074
rect 28590 55022 28642 55074
rect 30158 55022 30210 55074
rect 30494 55022 30546 55074
rect 31166 55022 31218 55074
rect 35534 55022 35586 55074
rect 42030 55022 42082 55074
rect 42142 55022 42194 55074
rect 42254 55022 42306 55074
rect 44942 55022 44994 55074
rect 45166 55022 45218 55074
rect 48078 55022 48130 55074
rect 51550 55022 51602 55074
rect 58158 55022 58210 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 27246 54686 27298 54738
rect 45054 54686 45106 54738
rect 47406 54686 47458 54738
rect 52334 54686 52386 54738
rect 1710 54574 1762 54626
rect 19406 54574 19458 54626
rect 21310 54574 21362 54626
rect 26350 54574 26402 54626
rect 29374 54574 29426 54626
rect 33182 54574 33234 54626
rect 34190 54574 34242 54626
rect 44718 54574 44770 54626
rect 44830 54574 44882 54626
rect 46846 54574 46898 54626
rect 49086 54574 49138 54626
rect 49310 54574 49362 54626
rect 50878 54574 50930 54626
rect 18622 54462 18674 54514
rect 20414 54462 20466 54514
rect 21198 54462 21250 54514
rect 22206 54462 22258 54514
rect 22430 54462 22482 54514
rect 23326 54462 23378 54514
rect 23662 54462 23714 54514
rect 25902 54462 25954 54514
rect 26798 54462 26850 54514
rect 27134 54462 27186 54514
rect 28142 54462 28194 54514
rect 28478 54462 28530 54514
rect 29038 54462 29090 54514
rect 30606 54462 30658 54514
rect 31950 54462 32002 54514
rect 34078 54462 34130 54514
rect 35646 54462 35698 54514
rect 37214 54462 37266 54514
rect 38110 54462 38162 54514
rect 41582 54462 41634 54514
rect 42254 54462 42306 54514
rect 43486 54462 43538 54514
rect 44382 54462 44434 54514
rect 46398 54462 46450 54514
rect 47070 54462 47122 54514
rect 47518 54462 47570 54514
rect 47630 54462 47682 54514
rect 49982 54462 50034 54514
rect 51550 54462 51602 54514
rect 19070 54350 19122 54402
rect 25678 54350 25730 54402
rect 27918 54350 27970 54402
rect 30158 54350 30210 54402
rect 35198 54350 35250 54402
rect 38446 54350 38498 54402
rect 41358 54350 41410 54402
rect 43822 54350 43874 54402
rect 46174 54350 46226 54402
rect 49198 54350 49250 54402
rect 50206 54350 50258 54402
rect 22094 54238 22146 54290
rect 22654 54238 22706 54290
rect 22766 54238 22818 54290
rect 23438 54238 23490 54290
rect 23774 54238 23826 54290
rect 25566 54238 25618 54290
rect 38670 54238 38722 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 41694 53902 41746 53954
rect 42254 53902 42306 53954
rect 42478 53902 42530 53954
rect 46174 53902 46226 53954
rect 47294 53902 47346 53954
rect 16830 53790 16882 53842
rect 19742 53790 19794 53842
rect 21422 53790 21474 53842
rect 23774 53790 23826 53842
rect 23886 53790 23938 53842
rect 28478 53790 28530 53842
rect 32958 53790 33010 53842
rect 34638 53790 34690 53842
rect 36094 53790 36146 53842
rect 37326 53790 37378 53842
rect 37998 53790 38050 53842
rect 39790 53790 39842 53842
rect 41358 53790 41410 53842
rect 46510 53790 46562 53842
rect 47854 53790 47906 53842
rect 50206 53790 50258 53842
rect 51326 53790 51378 53842
rect 16942 53678 16994 53730
rect 19294 53678 19346 53730
rect 19854 53678 19906 53730
rect 21758 53678 21810 53730
rect 22318 53678 22370 53730
rect 22542 53678 22594 53730
rect 22878 53678 22930 53730
rect 24782 53678 24834 53730
rect 25118 53678 25170 53730
rect 25790 53678 25842 53730
rect 26126 53678 26178 53730
rect 27918 53678 27970 53730
rect 29374 53678 29426 53730
rect 30046 53678 30098 53730
rect 30942 53678 30994 53730
rect 33294 53678 33346 53730
rect 33854 53678 33906 53730
rect 34414 53678 34466 53730
rect 34974 53678 35026 53730
rect 35870 53678 35922 53730
rect 37214 53678 37266 53730
rect 38782 53678 38834 53730
rect 39902 53678 39954 53730
rect 42030 53678 42082 53730
rect 42926 53678 42978 53730
rect 46958 53678 47010 53730
rect 47182 53678 47234 53730
rect 47966 53678 48018 53730
rect 49646 53678 49698 53730
rect 50094 53678 50146 53730
rect 50990 53678 51042 53730
rect 16046 53566 16098 53618
rect 16718 53566 16770 53618
rect 17838 53566 17890 53618
rect 23998 53566 24050 53618
rect 25454 53566 25506 53618
rect 27022 53566 27074 53618
rect 28366 53566 28418 53618
rect 29262 53566 29314 53618
rect 30270 53566 30322 53618
rect 33406 53566 33458 53618
rect 34190 53566 34242 53618
rect 39454 53566 39506 53618
rect 43598 53566 43650 53618
rect 43710 53566 43762 53618
rect 43934 53566 43986 53618
rect 48750 53566 48802 53618
rect 49086 53566 49138 53618
rect 49422 53566 49474 53618
rect 51662 53566 51714 53618
rect 52670 53566 52722 53618
rect 53006 53566 53058 53618
rect 16494 53454 16546 53506
rect 17166 53454 17218 53506
rect 17502 53454 17554 53506
rect 19406 53454 19458 53506
rect 19630 53454 19682 53506
rect 20414 53454 20466 53506
rect 20750 53454 20802 53506
rect 23102 53454 23154 53506
rect 25118 53454 25170 53506
rect 25902 53454 25954 53506
rect 26910 53454 26962 53506
rect 27694 53454 27746 53506
rect 28142 53454 28194 53506
rect 31502 53454 31554 53506
rect 36430 53454 36482 53506
rect 41582 53454 41634 53506
rect 46398 53454 46450 53506
rect 50318 53454 50370 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 20414 53118 20466 53170
rect 22766 53118 22818 53170
rect 23326 53118 23378 53170
rect 27806 53118 27858 53170
rect 28814 53118 28866 53170
rect 30830 53118 30882 53170
rect 33630 53118 33682 53170
rect 38894 53118 38946 53170
rect 39006 53118 39058 53170
rect 16606 53006 16658 53058
rect 17502 53006 17554 53058
rect 18622 53006 18674 53058
rect 18846 53006 18898 53058
rect 19630 53006 19682 53058
rect 20638 53006 20690 53058
rect 20750 53006 20802 53058
rect 28142 53006 28194 53058
rect 31278 53006 31330 53058
rect 38782 53006 38834 53058
rect 50654 53006 50706 53058
rect 58158 53006 58210 53058
rect 16718 52894 16770 52946
rect 17278 52894 17330 52946
rect 17614 52894 17666 52946
rect 18398 52894 18450 52946
rect 18510 52894 18562 52946
rect 19294 52894 19346 52946
rect 22094 52894 22146 52946
rect 22542 52894 22594 52946
rect 31054 52894 31106 52946
rect 31950 52894 32002 52946
rect 33406 52894 33458 52946
rect 33742 52894 33794 52946
rect 34190 52894 34242 52946
rect 34750 52894 34802 52946
rect 36766 52894 36818 52946
rect 47182 52894 47234 52946
rect 47406 52894 47458 52946
rect 50990 52894 51042 52946
rect 51774 52894 51826 52946
rect 21198 52782 21250 52834
rect 22318 52782 22370 52834
rect 22654 52782 22706 52834
rect 24558 52782 24610 52834
rect 26462 52782 26514 52834
rect 29262 52782 29314 52834
rect 30942 52782 30994 52834
rect 31726 52782 31778 52834
rect 32286 52782 32338 52834
rect 34638 52782 34690 52834
rect 36318 52782 36370 52834
rect 50878 52782 50930 52834
rect 51662 52782 51714 52834
rect 15598 52670 15650 52722
rect 15934 52670 15986 52722
rect 19182 52670 19234 52722
rect 19742 52670 19794 52722
rect 19966 52670 20018 52722
rect 20078 52670 20130 52722
rect 21870 52670 21922 52722
rect 35086 52670 35138 52722
rect 47630 52670 47682 52722
rect 48078 52670 48130 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 22990 52334 23042 52386
rect 23438 52334 23490 52386
rect 31278 52334 31330 52386
rect 43598 52334 43650 52386
rect 47966 52334 48018 52386
rect 15822 52222 15874 52274
rect 19070 52222 19122 52274
rect 19630 52222 19682 52274
rect 21422 52222 21474 52274
rect 25342 52222 25394 52274
rect 27470 52222 27522 52274
rect 34190 52222 34242 52274
rect 40014 52222 40066 52274
rect 40910 52222 40962 52274
rect 43262 52222 43314 52274
rect 51326 52222 51378 52274
rect 51774 52222 51826 52274
rect 16382 52110 16434 52162
rect 16942 52110 16994 52162
rect 19406 52110 19458 52162
rect 20862 52110 20914 52162
rect 21870 52110 21922 52162
rect 22094 52110 22146 52162
rect 22766 52110 22818 52162
rect 23662 52110 23714 52162
rect 23998 52110 24050 52162
rect 24558 52110 24610 52162
rect 25566 52110 25618 52162
rect 26910 52110 26962 52162
rect 27694 52110 27746 52162
rect 20526 51998 20578 52050
rect 20638 51998 20690 52050
rect 25006 51998 25058 52050
rect 25342 51998 25394 52050
rect 27134 51998 27186 52050
rect 28366 51998 28418 52050
rect 28702 52110 28754 52162
rect 30494 52110 30546 52162
rect 34078 52110 34130 52162
rect 34302 52110 34354 52162
rect 34638 52110 34690 52162
rect 38446 52110 38498 52162
rect 39118 52110 39170 52162
rect 40574 52110 40626 52162
rect 42030 52110 42082 52162
rect 42254 52110 42306 52162
rect 43150 52110 43202 52162
rect 43486 52110 43538 52162
rect 51438 52110 51490 52162
rect 31166 51998 31218 52050
rect 31278 51998 31330 52050
rect 38558 51998 38610 52050
rect 45726 51998 45778 52050
rect 47630 51998 47682 52050
rect 47854 51998 47906 52050
rect 15486 51886 15538 51938
rect 15710 51886 15762 51938
rect 15934 51886 15986 51938
rect 23886 51886 23938 51938
rect 24110 51886 24162 51938
rect 27246 51886 27298 51938
rect 29262 51886 29314 51938
rect 30830 51886 30882 51938
rect 39454 51886 39506 51938
rect 39902 51886 39954 51938
rect 40126 51886 40178 51938
rect 40798 51886 40850 51938
rect 41022 51886 41074 51938
rect 41246 51886 41298 51938
rect 45838 51886 45890 51938
rect 46062 51886 46114 51938
rect 50990 51886 51042 51938
rect 51214 51886 51266 51938
rect 51886 51886 51938 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 22990 51550 23042 51602
rect 23886 51550 23938 51602
rect 24558 51550 24610 51602
rect 25678 51550 25730 51602
rect 39454 51550 39506 51602
rect 41022 51550 41074 51602
rect 47294 51550 47346 51602
rect 51662 51550 51714 51602
rect 16494 51438 16546 51490
rect 19182 51438 19234 51490
rect 23214 51438 23266 51490
rect 23662 51438 23714 51490
rect 28366 51438 28418 51490
rect 28478 51438 28530 51490
rect 36990 51438 37042 51490
rect 37550 51438 37602 51490
rect 38334 51438 38386 51490
rect 38782 51438 38834 51490
rect 41134 51438 41186 51490
rect 42702 51438 42754 51490
rect 46174 51438 46226 51490
rect 47406 51438 47458 51490
rect 51102 51438 51154 51490
rect 53902 51438 53954 51490
rect 58158 51438 58210 51490
rect 15150 51326 15202 51378
rect 15486 51326 15538 51378
rect 15934 51326 15986 51378
rect 16270 51326 16322 51378
rect 16718 51326 16770 51378
rect 19070 51326 19122 51378
rect 20974 51326 21026 51378
rect 22542 51326 22594 51378
rect 24110 51326 24162 51378
rect 25118 51326 25170 51378
rect 25566 51326 25618 51378
rect 25790 51326 25842 51378
rect 26462 51326 26514 51378
rect 27246 51326 27298 51378
rect 27806 51326 27858 51378
rect 28142 51326 28194 51378
rect 28926 51326 28978 51378
rect 29262 51326 29314 51378
rect 30606 51326 30658 51378
rect 30830 51326 30882 51378
rect 31054 51326 31106 51378
rect 31278 51326 31330 51378
rect 34302 51326 34354 51378
rect 36094 51326 36146 51378
rect 36430 51326 36482 51378
rect 37886 51326 37938 51378
rect 39118 51326 39170 51378
rect 42030 51326 42082 51378
rect 43374 51326 43426 51378
rect 45726 51326 45778 51378
rect 46958 51326 47010 51378
rect 47070 51326 47122 51378
rect 50878 51326 50930 51378
rect 51550 51326 51602 51378
rect 52782 51326 52834 51378
rect 53230 51326 53282 51378
rect 53566 51326 53618 51378
rect 15598 51214 15650 51266
rect 16382 51214 16434 51266
rect 17502 51214 17554 51266
rect 18398 51214 18450 51266
rect 18734 51214 18786 51266
rect 23998 51214 24050 51266
rect 26910 51214 26962 51266
rect 28254 51214 28306 51266
rect 29822 51214 29874 51266
rect 31166 51214 31218 51266
rect 34078 51214 34130 51266
rect 42254 51214 42306 51266
rect 43262 51214 43314 51266
rect 44046 51214 44098 51266
rect 45502 51214 45554 51266
rect 52334 51214 52386 51266
rect 24334 51102 24386 51154
rect 24782 51102 24834 51154
rect 34750 51102 34802 51154
rect 37886 51102 37938 51154
rect 40910 51102 40962 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 15486 50766 15538 50818
rect 16382 50766 16434 50818
rect 17726 50766 17778 50818
rect 18062 50766 18114 50818
rect 19518 50766 19570 50818
rect 25342 50766 25394 50818
rect 34862 50766 34914 50818
rect 42142 50766 42194 50818
rect 42478 50766 42530 50818
rect 47406 50766 47458 50818
rect 52782 50766 52834 50818
rect 57934 50766 57986 50818
rect 12910 50654 12962 50706
rect 15150 50654 15202 50706
rect 17390 50654 17442 50706
rect 20190 50654 20242 50706
rect 22542 50654 22594 50706
rect 23886 50654 23938 50706
rect 27582 50654 27634 50706
rect 39230 50654 39282 50706
rect 44942 50654 44994 50706
rect 13470 50542 13522 50594
rect 14142 50542 14194 50594
rect 18846 50542 18898 50594
rect 22094 50542 22146 50594
rect 22318 50542 22370 50594
rect 25230 50542 25282 50594
rect 25566 50542 25618 50594
rect 29150 50542 29202 50594
rect 29486 50542 29538 50594
rect 31166 50542 31218 50594
rect 33294 50542 33346 50594
rect 33966 50542 34018 50594
rect 34526 50542 34578 50594
rect 38782 50542 38834 50594
rect 39342 50542 39394 50594
rect 42478 50542 42530 50594
rect 44046 50542 44098 50594
rect 45166 50542 45218 50594
rect 46622 50542 46674 50594
rect 46846 50542 46898 50594
rect 47742 50542 47794 50594
rect 48638 50542 48690 50594
rect 50430 50542 50482 50594
rect 51662 50542 51714 50594
rect 52894 50542 52946 50594
rect 55582 50542 55634 50594
rect 14590 50430 14642 50482
rect 14814 50430 14866 50482
rect 15038 50430 15090 50482
rect 15262 50430 15314 50482
rect 16942 50430 16994 50482
rect 18622 50430 18674 50482
rect 19406 50430 19458 50482
rect 19518 50430 19570 50482
rect 20526 50430 20578 50482
rect 20638 50430 20690 50482
rect 20862 50430 20914 50482
rect 22654 50430 22706 50482
rect 22990 50430 23042 50482
rect 23102 50430 23154 50482
rect 23774 50430 23826 50482
rect 25006 50430 25058 50482
rect 26462 50430 26514 50482
rect 27694 50430 27746 50482
rect 28142 50430 28194 50482
rect 30382 50430 30434 50482
rect 31054 50430 31106 50482
rect 31502 50430 31554 50482
rect 31726 50430 31778 50482
rect 31838 50430 31890 50482
rect 32958 50430 33010 50482
rect 33070 50430 33122 50482
rect 33854 50430 33906 50482
rect 39006 50430 39058 50482
rect 39902 50430 39954 50482
rect 44158 50430 44210 50482
rect 44382 50430 44434 50482
rect 45838 50430 45890 50482
rect 46958 50430 47010 50482
rect 48078 50430 48130 50482
rect 50766 50430 50818 50482
rect 51102 50430 51154 50482
rect 52782 50430 52834 50482
rect 13582 50318 13634 50370
rect 13694 50318 13746 50370
rect 15710 50318 15762 50370
rect 16382 50318 16434 50370
rect 16606 50318 16658 50370
rect 17950 50318 18002 50370
rect 18958 50318 19010 50370
rect 19182 50318 19234 50370
rect 21422 50318 21474 50370
rect 23326 50318 23378 50370
rect 23998 50318 24050 50370
rect 28702 50318 28754 50370
rect 29598 50318 29650 50370
rect 29710 50318 29762 50370
rect 48638 50318 48690 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 19294 49982 19346 50034
rect 21086 49982 21138 50034
rect 27022 49982 27074 50034
rect 29822 49982 29874 50034
rect 30606 49982 30658 50034
rect 34190 49982 34242 50034
rect 35422 49982 35474 50034
rect 38110 49982 38162 50034
rect 47518 49982 47570 50034
rect 50430 49982 50482 50034
rect 12462 49870 12514 49922
rect 16270 49870 16322 49922
rect 16382 49870 16434 49922
rect 17838 49870 17890 49922
rect 18398 49870 18450 49922
rect 19630 49870 19682 49922
rect 20414 49870 20466 49922
rect 21198 49870 21250 49922
rect 24110 49870 24162 49922
rect 25342 49870 25394 49922
rect 30046 49870 30098 49922
rect 35534 49870 35586 49922
rect 36878 49870 36930 49922
rect 39902 49870 39954 49922
rect 43038 49870 43090 49922
rect 43150 49870 43202 49922
rect 45054 49870 45106 49922
rect 46846 49870 46898 49922
rect 47854 49870 47906 49922
rect 58158 49870 58210 49922
rect 13134 49758 13186 49810
rect 13806 49758 13858 49810
rect 16046 49758 16098 49810
rect 16718 49758 16770 49810
rect 17502 49758 17554 49810
rect 18958 49758 19010 49810
rect 19406 49758 19458 49810
rect 20190 49758 20242 49810
rect 21422 49758 21474 49810
rect 21870 49758 21922 49810
rect 22430 49758 22482 49810
rect 23214 49758 23266 49810
rect 25230 49758 25282 49810
rect 26126 49758 26178 49810
rect 26686 49758 26738 49810
rect 28030 49758 28082 49810
rect 29598 49758 29650 49810
rect 30270 49758 30322 49810
rect 30718 49758 30770 49810
rect 30830 49758 30882 49810
rect 31166 49758 31218 49810
rect 34414 49758 34466 49810
rect 35758 49758 35810 49810
rect 36542 49758 36594 49810
rect 37438 49758 37490 49810
rect 37886 49758 37938 49810
rect 39566 49758 39618 49810
rect 43374 49758 43426 49810
rect 45390 49758 45442 49810
rect 45950 49758 46002 49810
rect 47182 49758 47234 49810
rect 47630 49758 47682 49810
rect 49870 49758 49922 49810
rect 11230 49646 11282 49698
rect 11678 49646 11730 49698
rect 12126 49646 12178 49698
rect 13470 49646 13522 49698
rect 14702 49646 14754 49698
rect 15710 49646 15762 49698
rect 16830 49646 16882 49698
rect 23550 49646 23602 49698
rect 24222 49646 24274 49698
rect 24670 49646 24722 49698
rect 25454 49646 25506 49698
rect 28590 49646 28642 49698
rect 29262 49646 29314 49698
rect 30046 49646 30098 49698
rect 36430 49646 36482 49698
rect 37998 49646 38050 49698
rect 46062 49646 46114 49698
rect 50094 49646 50146 49698
rect 11118 49534 11170 49586
rect 11678 49534 11730 49586
rect 12014 49534 12066 49586
rect 12350 49534 12402 49586
rect 14030 49534 14082 49586
rect 22990 49534 23042 49586
rect 23886 49534 23938 49586
rect 34078 49534 34130 49586
rect 35422 49534 35474 49586
rect 45390 49534 45442 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 19742 49198 19794 49250
rect 35870 49198 35922 49250
rect 44270 49198 44322 49250
rect 47854 49198 47906 49250
rect 49758 49198 49810 49250
rect 50990 49198 51042 49250
rect 13582 49086 13634 49138
rect 14590 49086 14642 49138
rect 17838 49086 17890 49138
rect 19294 49086 19346 49138
rect 20750 49086 20802 49138
rect 21758 49086 21810 49138
rect 29262 49086 29314 49138
rect 39006 49086 39058 49138
rect 39566 49086 39618 49138
rect 40238 49086 40290 49138
rect 43598 49086 43650 49138
rect 48974 49086 49026 49138
rect 50094 49086 50146 49138
rect 58158 49086 58210 49138
rect 16158 48974 16210 49026
rect 16606 48974 16658 49026
rect 17166 48974 17218 49026
rect 18958 48974 19010 49026
rect 21310 48974 21362 49026
rect 21646 48974 21698 49026
rect 21870 48974 21922 49026
rect 23774 48974 23826 49026
rect 25454 48974 25506 49026
rect 26238 48974 26290 49026
rect 27358 48974 27410 49026
rect 30046 48974 30098 49026
rect 30830 48974 30882 49026
rect 31278 48974 31330 49026
rect 33182 48974 33234 49026
rect 33406 48974 33458 49026
rect 33630 48974 33682 49026
rect 34078 48974 34130 49026
rect 34526 48974 34578 49026
rect 34974 48974 35026 49026
rect 35422 48974 35474 49026
rect 35758 48974 35810 49026
rect 39454 48974 39506 49026
rect 42254 48974 42306 49026
rect 42814 48974 42866 49026
rect 43262 48974 43314 49026
rect 45950 48974 46002 49026
rect 46174 48974 46226 49026
rect 46510 48974 46562 49026
rect 49870 48974 49922 49026
rect 22542 48862 22594 48914
rect 22878 48862 22930 48914
rect 23550 48862 23602 48914
rect 26462 48862 26514 48914
rect 30270 48862 30322 48914
rect 42926 48862 42978 48914
rect 43934 48862 43986 48914
rect 47518 48862 47570 48914
rect 47742 48862 47794 48914
rect 49086 48862 49138 48914
rect 50878 48862 50930 48914
rect 14030 48750 14082 48802
rect 22206 48750 22258 48802
rect 23214 48750 23266 48802
rect 27134 48750 27186 48802
rect 28030 48750 28082 48802
rect 28590 48750 28642 48802
rect 29710 48750 29762 48802
rect 31390 48750 31442 48802
rect 33294 48750 33346 48802
rect 37774 48750 37826 48802
rect 43486 48750 43538 48802
rect 44158 48750 44210 48802
rect 46062 48750 46114 48802
rect 50990 48750 51042 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 21646 48414 21698 48466
rect 23326 48414 23378 48466
rect 25790 48414 25842 48466
rect 32174 48414 32226 48466
rect 34190 48414 34242 48466
rect 35646 48414 35698 48466
rect 35870 48414 35922 48466
rect 38446 48414 38498 48466
rect 39678 48414 39730 48466
rect 42366 48414 42418 48466
rect 44942 48414 44994 48466
rect 20190 48302 20242 48354
rect 22654 48302 22706 48354
rect 25902 48302 25954 48354
rect 27246 48302 27298 48354
rect 29934 48302 29986 48354
rect 30158 48302 30210 48354
rect 30494 48302 30546 48354
rect 31278 48302 31330 48354
rect 34078 48302 34130 48354
rect 35534 48302 35586 48354
rect 36430 48302 36482 48354
rect 37998 48302 38050 48354
rect 38558 48302 38610 48354
rect 40014 48302 40066 48354
rect 42142 48302 42194 48354
rect 42478 48302 42530 48354
rect 44046 48302 44098 48354
rect 45614 48302 45666 48354
rect 11230 48190 11282 48242
rect 11678 48190 11730 48242
rect 13358 48190 13410 48242
rect 13806 48190 13858 48242
rect 14142 48190 14194 48242
rect 15374 48190 15426 48242
rect 20414 48190 20466 48242
rect 21534 48190 21586 48242
rect 26462 48190 26514 48242
rect 27470 48190 27522 48242
rect 28142 48190 28194 48242
rect 28926 48190 28978 48242
rect 29486 48190 29538 48242
rect 30830 48190 30882 48242
rect 31166 48190 31218 48242
rect 32062 48190 32114 48242
rect 36318 48190 36370 48242
rect 36542 48190 36594 48242
rect 37214 48190 37266 48242
rect 38334 48190 38386 48242
rect 38894 48190 38946 48242
rect 39118 48190 39170 48242
rect 39454 48190 39506 48242
rect 40238 48190 40290 48242
rect 42590 48190 42642 48242
rect 43934 48190 43986 48242
rect 44942 48190 44994 48242
rect 49758 48190 49810 48242
rect 49982 48190 50034 48242
rect 15486 48078 15538 48130
rect 16270 48078 16322 48130
rect 18510 48078 18562 48130
rect 19294 48078 19346 48130
rect 24110 48078 24162 48130
rect 24782 48078 24834 48130
rect 25342 48078 25394 48130
rect 26910 48078 26962 48130
rect 41022 48078 41074 48130
rect 45726 48078 45778 48130
rect 50654 48078 50706 48130
rect 23214 47966 23266 48018
rect 23550 47966 23602 48018
rect 25678 47966 25730 48018
rect 28926 47966 28978 48018
rect 29822 47966 29874 48018
rect 34302 47966 34354 48018
rect 39342 47966 39394 48018
rect 45390 47966 45442 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 16606 47630 16658 47682
rect 25342 47630 25394 47682
rect 26798 47630 26850 47682
rect 30158 47630 30210 47682
rect 30942 47630 30994 47682
rect 13918 47518 13970 47570
rect 16718 47518 16770 47570
rect 17614 47518 17666 47570
rect 19630 47518 19682 47570
rect 22318 47518 22370 47570
rect 22990 47518 23042 47570
rect 24334 47518 24386 47570
rect 31614 47630 31666 47682
rect 39790 47630 39842 47682
rect 27358 47518 27410 47570
rect 29934 47518 29986 47570
rect 31390 47518 31442 47570
rect 31950 47518 32002 47570
rect 37438 47518 37490 47570
rect 49310 47518 49362 47570
rect 50430 47518 50482 47570
rect 57934 47518 57986 47570
rect 13582 47406 13634 47458
rect 16270 47406 16322 47458
rect 17278 47406 17330 47458
rect 18734 47406 18786 47458
rect 19070 47406 19122 47458
rect 21534 47406 21586 47458
rect 23998 47406 24050 47458
rect 24446 47406 24498 47458
rect 24782 47406 24834 47458
rect 27022 47406 27074 47458
rect 27470 47406 27522 47458
rect 27582 47406 27634 47458
rect 28142 47406 28194 47458
rect 29262 47406 29314 47458
rect 30270 47406 30322 47458
rect 32062 47406 32114 47458
rect 36542 47406 36594 47458
rect 37214 47406 37266 47458
rect 39566 47406 39618 47458
rect 39902 47406 39954 47458
rect 46622 47406 46674 47458
rect 49534 47406 49586 47458
rect 50654 47406 50706 47458
rect 55582 47406 55634 47458
rect 18510 47294 18562 47346
rect 19742 47294 19794 47346
rect 20526 47294 20578 47346
rect 20638 47294 20690 47346
rect 23550 47294 23602 47346
rect 24222 47294 24274 47346
rect 27246 47294 27298 47346
rect 28254 47294 28306 47346
rect 36206 47294 36258 47346
rect 38110 47294 38162 47346
rect 39342 47294 39394 47346
rect 45502 47294 45554 47346
rect 46958 47294 47010 47346
rect 51326 47294 51378 47346
rect 12350 47182 12402 47234
rect 13022 47182 13074 47234
rect 14702 47182 14754 47234
rect 15598 47182 15650 47234
rect 18174 47182 18226 47234
rect 19518 47182 19570 47234
rect 20302 47182 20354 47234
rect 22766 47182 22818 47234
rect 22878 47182 22930 47234
rect 23326 47182 23378 47234
rect 23438 47182 23490 47234
rect 25342 47182 25394 47234
rect 25678 47182 25730 47234
rect 26126 47182 26178 47234
rect 26686 47182 26738 47234
rect 28030 47182 28082 47234
rect 28478 47182 28530 47234
rect 31166 47182 31218 47234
rect 36318 47182 36370 47234
rect 40126 47182 40178 47234
rect 45614 47182 45666 47234
rect 46846 47182 46898 47234
rect 49870 47182 49922 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 16046 46846 16098 46898
rect 16830 46846 16882 46898
rect 19070 46846 19122 46898
rect 23774 46846 23826 46898
rect 24222 46846 24274 46898
rect 25342 46846 25394 46898
rect 31278 46846 31330 46898
rect 31390 46846 31442 46898
rect 35422 46846 35474 46898
rect 41022 46846 41074 46898
rect 14030 46734 14082 46786
rect 14366 46734 14418 46786
rect 15038 46734 15090 46786
rect 18062 46734 18114 46786
rect 18846 46734 18898 46786
rect 20974 46734 21026 46786
rect 21310 46734 21362 46786
rect 21422 46734 21474 46786
rect 23102 46734 23154 46786
rect 23662 46734 23714 46786
rect 23886 46734 23938 46786
rect 24446 46734 24498 46786
rect 24558 46734 24610 46786
rect 35086 46734 35138 46786
rect 42030 46734 42082 46786
rect 42926 46734 42978 46786
rect 44158 46734 44210 46786
rect 45166 46734 45218 46786
rect 46510 46734 46562 46786
rect 51102 46734 51154 46786
rect 52446 46734 52498 46786
rect 11678 46622 11730 46674
rect 13022 46622 13074 46674
rect 13806 46622 13858 46674
rect 14702 46622 14754 46674
rect 17726 46622 17778 46674
rect 17838 46622 17890 46674
rect 19406 46622 19458 46674
rect 19854 46622 19906 46674
rect 20638 46622 20690 46674
rect 21646 46622 21698 46674
rect 21870 46622 21922 46674
rect 22542 46622 22594 46674
rect 27246 46622 27298 46674
rect 27694 46622 27746 46674
rect 30830 46622 30882 46674
rect 31166 46622 31218 46674
rect 41358 46622 41410 46674
rect 41806 46622 41858 46674
rect 42590 46622 42642 46674
rect 43150 46622 43202 46674
rect 43934 46622 43986 46674
rect 45054 46622 45106 46674
rect 45390 46622 45442 46674
rect 47518 46622 47570 46674
rect 50654 46622 50706 46674
rect 51326 46622 51378 46674
rect 51438 46622 51490 46674
rect 52894 46622 52946 46674
rect 53342 46622 53394 46674
rect 11230 46510 11282 46562
rect 12350 46510 12402 46562
rect 15486 46510 15538 46562
rect 16270 46510 16322 46562
rect 17950 46510 18002 46562
rect 20302 46510 20354 46562
rect 22654 46510 22706 46562
rect 25790 46510 25842 46562
rect 26686 46510 26738 46562
rect 28142 46510 28194 46562
rect 28702 46510 28754 46562
rect 29038 46510 29090 46562
rect 30494 46510 30546 46562
rect 42142 46510 42194 46562
rect 44606 46510 44658 46562
rect 46062 46510 46114 46562
rect 48190 46510 48242 46562
rect 53118 46510 53170 46562
rect 12686 46398 12738 46450
rect 13022 46398 13074 46450
rect 16494 46398 16546 46450
rect 17390 46398 17442 46450
rect 19182 46398 19234 46450
rect 27022 46398 27074 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 13694 46062 13746 46114
rect 18622 46062 18674 46114
rect 19966 46062 20018 46114
rect 32734 46062 32786 46114
rect 35870 46062 35922 46114
rect 51662 46062 51714 46114
rect 11902 45950 11954 46002
rect 12462 45950 12514 46002
rect 16046 45950 16098 46002
rect 18286 45950 18338 46002
rect 35198 45950 35250 46002
rect 11566 45838 11618 45890
rect 13470 45838 13522 45890
rect 14030 45838 14082 45890
rect 14142 45838 14194 45890
rect 14254 45838 14306 45890
rect 14366 45838 14418 45890
rect 14926 45838 14978 45890
rect 15486 45838 15538 45890
rect 16270 45838 16322 45890
rect 16606 45838 16658 45890
rect 16942 45838 16994 45890
rect 17390 45838 17442 45890
rect 17502 45838 17554 45890
rect 17614 45838 17666 45890
rect 17726 45838 17778 45890
rect 17950 45838 18002 45890
rect 19742 45838 19794 45890
rect 20078 45838 20130 45890
rect 21870 45838 21922 45890
rect 23102 45838 23154 45890
rect 23438 45838 23490 45890
rect 23774 45838 23826 45890
rect 26686 45838 26738 45890
rect 27022 45838 27074 45890
rect 27470 45838 27522 45890
rect 28366 45838 28418 45890
rect 31166 45838 31218 45890
rect 31614 45838 31666 45890
rect 32510 45838 32562 45890
rect 32846 45838 32898 45890
rect 33518 45838 33570 45890
rect 35086 45838 35138 45890
rect 39118 45838 39170 45890
rect 43822 45838 43874 45890
rect 44046 45838 44098 45890
rect 45390 45838 45442 45890
rect 45726 45838 45778 45890
rect 46510 45838 46562 45890
rect 46846 45838 46898 45890
rect 47070 45838 47122 45890
rect 49534 45838 49586 45890
rect 49870 45838 49922 45890
rect 50318 45838 50370 45890
rect 51662 45838 51714 45890
rect 52894 45838 52946 45890
rect 16718 45726 16770 45778
rect 18510 45726 18562 45778
rect 25230 45726 25282 45778
rect 27694 45726 27746 45778
rect 27806 45726 27858 45778
rect 28030 45726 28082 45778
rect 29262 45726 29314 45778
rect 30046 45726 30098 45778
rect 30942 45726 30994 45778
rect 31838 45726 31890 45778
rect 33742 45726 33794 45778
rect 34302 45726 34354 45778
rect 38558 45726 38610 45778
rect 38894 45726 38946 45778
rect 39454 45726 39506 45778
rect 43710 45726 43762 45778
rect 44270 45726 44322 45778
rect 45502 45726 45554 45778
rect 51326 45726 51378 45778
rect 53118 45726 53170 45778
rect 12910 45614 12962 45666
rect 19070 45614 19122 45666
rect 19518 45614 19570 45666
rect 20302 45614 20354 45666
rect 20750 45614 20802 45666
rect 26686 45614 26738 45666
rect 27246 45614 27298 45666
rect 28142 45614 28194 45666
rect 29710 45614 29762 45666
rect 30606 45614 30658 45666
rect 33966 45614 34018 45666
rect 40126 45614 40178 45666
rect 40462 45614 40514 45666
rect 46734 45614 46786 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 10558 45278 10610 45330
rect 17390 45278 17442 45330
rect 18398 45278 18450 45330
rect 18846 45278 18898 45330
rect 26462 45278 26514 45330
rect 26686 45278 26738 45330
rect 28030 45278 28082 45330
rect 31726 45278 31778 45330
rect 34638 45278 34690 45330
rect 40014 45278 40066 45330
rect 42702 45278 42754 45330
rect 44830 45278 44882 45330
rect 10894 45166 10946 45218
rect 16718 45166 16770 45218
rect 19966 45166 20018 45218
rect 24446 45166 24498 45218
rect 25342 45166 25394 45218
rect 26014 45166 26066 45218
rect 29038 45166 29090 45218
rect 30046 45166 30098 45218
rect 30830 45166 30882 45218
rect 37998 45166 38050 45218
rect 41918 45166 41970 45218
rect 46398 45166 46450 45218
rect 11342 45054 11394 45106
rect 11902 45054 11954 45106
rect 13022 45054 13074 45106
rect 14366 45054 14418 45106
rect 15038 45054 15090 45106
rect 16270 45054 16322 45106
rect 19854 45054 19906 45106
rect 20190 45054 20242 45106
rect 22766 45054 22818 45106
rect 23886 45054 23938 45106
rect 24334 45054 24386 45106
rect 25678 45054 25730 45106
rect 27022 45054 27074 45106
rect 27470 45054 27522 45106
rect 27806 45054 27858 45106
rect 28590 45054 28642 45106
rect 29486 45054 29538 45106
rect 30606 45054 30658 45106
rect 34190 45054 34242 45106
rect 34414 45054 34466 45106
rect 34862 45054 34914 45106
rect 37886 45054 37938 45106
rect 38222 45054 38274 45106
rect 38558 45054 38610 45106
rect 38782 45054 38834 45106
rect 39454 45054 39506 45106
rect 39790 45054 39842 45106
rect 41246 45054 41298 45106
rect 42254 45054 42306 45106
rect 42478 45054 42530 45106
rect 44606 45054 44658 45106
rect 46286 45054 46338 45106
rect 46622 45054 46674 45106
rect 49758 45054 49810 45106
rect 11118 44942 11170 44994
rect 14478 44942 14530 44994
rect 17838 44942 17890 44994
rect 22094 44942 22146 44994
rect 22654 44942 22706 44994
rect 26798 44942 26850 44994
rect 32286 44942 32338 44994
rect 35198 44942 35250 44994
rect 41022 44942 41074 44994
rect 42366 44942 42418 44994
rect 49534 44942 49586 44994
rect 23662 44830 23714 44882
rect 24446 44830 24498 44882
rect 28142 44830 28194 44882
rect 29710 44830 29762 44882
rect 31390 44830 31442 44882
rect 40126 44830 40178 44882
rect 50094 44830 50146 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 15822 44494 15874 44546
rect 37326 44494 37378 44546
rect 50878 44494 50930 44546
rect 12238 44382 12290 44434
rect 14366 44382 14418 44434
rect 22430 44382 22482 44434
rect 29262 44382 29314 44434
rect 34862 44382 34914 44434
rect 39118 44382 39170 44434
rect 39678 44382 39730 44434
rect 42702 44382 42754 44434
rect 46174 44382 46226 44434
rect 47518 44382 47570 44434
rect 57934 44382 57986 44434
rect 10110 44270 10162 44322
rect 10894 44270 10946 44322
rect 14590 44270 14642 44322
rect 14926 44270 14978 44322
rect 15150 44270 15202 44322
rect 15934 44270 15986 44322
rect 16942 44270 16994 44322
rect 20750 44270 20802 44322
rect 21310 44270 21362 44322
rect 21758 44270 21810 44322
rect 23662 44270 23714 44322
rect 25006 44270 25058 44322
rect 25342 44270 25394 44322
rect 26574 44270 26626 44322
rect 28254 44270 28306 44322
rect 29822 44270 29874 44322
rect 31166 44270 31218 44322
rect 31502 44270 31554 44322
rect 34638 44270 34690 44322
rect 35310 44270 35362 44322
rect 36990 44270 37042 44322
rect 37326 44270 37378 44322
rect 38670 44270 38722 44322
rect 42366 44270 42418 44322
rect 43486 44270 43538 44322
rect 45950 44270 46002 44322
rect 46846 44270 46898 44322
rect 47406 44270 47458 44322
rect 51214 44270 51266 44322
rect 55582 44270 55634 44322
rect 10782 44158 10834 44210
rect 17054 44158 17106 44210
rect 19630 44158 19682 44210
rect 22094 44158 22146 44210
rect 27134 44158 27186 44210
rect 31838 44158 31890 44210
rect 39230 44158 39282 44210
rect 42702 44158 42754 44210
rect 48302 44158 48354 44210
rect 52670 44158 52722 44210
rect 53006 44158 53058 44210
rect 10334 44046 10386 44098
rect 14702 44046 14754 44098
rect 15486 44046 15538 44098
rect 15710 44046 15762 44098
rect 16382 44046 16434 44098
rect 16494 44046 16546 44098
rect 16606 44046 16658 44098
rect 20526 44046 20578 44098
rect 22990 44046 23042 44098
rect 26910 44046 26962 44098
rect 38334 44046 38386 44098
rect 39006 44046 39058 44098
rect 50990 44046 51042 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 18846 43710 18898 43762
rect 31278 43710 31330 43762
rect 43038 43710 43090 43762
rect 47406 43710 47458 43762
rect 47630 43710 47682 43762
rect 50542 43710 50594 43762
rect 12462 43598 12514 43650
rect 13582 43598 13634 43650
rect 13694 43598 13746 43650
rect 16382 43598 16434 43650
rect 16830 43598 16882 43650
rect 17502 43598 17554 43650
rect 17614 43598 17666 43650
rect 19070 43598 19122 43650
rect 27246 43598 27298 43650
rect 27470 43598 27522 43650
rect 28590 43598 28642 43650
rect 29710 43598 29762 43650
rect 33854 43598 33906 43650
rect 34750 43598 34802 43650
rect 35758 43598 35810 43650
rect 38782 43598 38834 43650
rect 41022 43598 41074 43650
rect 42814 43598 42866 43650
rect 49758 43598 49810 43650
rect 50654 43598 50706 43650
rect 10222 43486 10274 43538
rect 10446 43486 10498 43538
rect 10894 43486 10946 43538
rect 11566 43486 11618 43538
rect 12126 43486 12178 43538
rect 15710 43486 15762 43538
rect 17726 43486 17778 43538
rect 18734 43486 18786 43538
rect 19518 43486 19570 43538
rect 20526 43486 20578 43538
rect 22206 43486 22258 43538
rect 23550 43486 23602 43538
rect 25230 43486 25282 43538
rect 26798 43486 26850 43538
rect 27582 43486 27634 43538
rect 29150 43486 29202 43538
rect 30270 43486 30322 43538
rect 30718 43486 30770 43538
rect 31054 43486 31106 43538
rect 32286 43486 32338 43538
rect 34302 43486 34354 43538
rect 35870 43486 35922 43538
rect 38110 43486 38162 43538
rect 42030 43486 42082 43538
rect 44942 43486 44994 43538
rect 47070 43486 47122 43538
rect 47518 43486 47570 43538
rect 50430 43486 50482 43538
rect 51214 43486 51266 43538
rect 52334 43486 52386 43538
rect 11902 43374 11954 43426
rect 13022 43374 13074 43426
rect 14590 43374 14642 43426
rect 18398 43374 18450 43426
rect 19294 43374 19346 43426
rect 20302 43374 20354 43426
rect 23886 43374 23938 43426
rect 25566 43374 25618 43426
rect 28142 43374 28194 43426
rect 31950 43374 32002 43426
rect 36206 43374 36258 43426
rect 37886 43374 37938 43426
rect 39230 43374 39282 43426
rect 41582 43374 41634 43426
rect 42366 43374 42418 43426
rect 45166 43374 45218 43426
rect 50990 43374 51042 43426
rect 52446 43374 52498 43426
rect 10894 43262 10946 43314
rect 11006 43262 11058 43314
rect 13694 43262 13746 43314
rect 19854 43262 19906 43314
rect 21758 43262 21810 43314
rect 25454 43262 25506 43314
rect 26910 43262 26962 43314
rect 43150 43262 43202 43314
rect 45278 43262 45330 43314
rect 49534 43262 49586 43314
rect 49870 43262 49922 43314
rect 52670 43262 52722 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 15038 42926 15090 42978
rect 17390 42926 17442 42978
rect 18846 42926 18898 42978
rect 29374 42926 29426 42978
rect 29710 42926 29762 42978
rect 10110 42814 10162 42866
rect 11230 42814 11282 42866
rect 15598 42814 15650 42866
rect 16606 42814 16658 42866
rect 21646 42814 21698 42866
rect 22542 42814 22594 42866
rect 23438 42814 23490 42866
rect 24558 42814 24610 42866
rect 25790 42814 25842 42866
rect 26574 42814 26626 42866
rect 27022 42814 27074 42866
rect 28142 42814 28194 42866
rect 30830 42814 30882 42866
rect 31726 42814 31778 42866
rect 32622 42814 32674 42866
rect 34302 42814 34354 42866
rect 35198 42814 35250 42866
rect 37550 42814 37602 42866
rect 38110 42814 38162 42866
rect 41806 42814 41858 42866
rect 43150 42814 43202 42866
rect 57934 42814 57986 42866
rect 10446 42702 10498 42754
rect 13470 42702 13522 42754
rect 15710 42702 15762 42754
rect 18174 42702 18226 42754
rect 18958 42702 19010 42754
rect 19630 42702 19682 42754
rect 19854 42702 19906 42754
rect 20302 42702 20354 42754
rect 21758 42702 21810 42754
rect 21982 42702 22034 42754
rect 24670 42702 24722 42754
rect 30606 42702 30658 42754
rect 34974 42702 35026 42754
rect 36318 42702 36370 42754
rect 38446 42702 38498 42754
rect 38558 42702 38610 42754
rect 39006 42702 39058 42754
rect 39454 42702 39506 42754
rect 39902 42702 39954 42754
rect 40014 42702 40066 42754
rect 40238 42702 40290 42754
rect 42030 42702 42082 42754
rect 45390 42702 45442 42754
rect 45502 42702 45554 42754
rect 46174 42702 46226 42754
rect 49198 42702 49250 42754
rect 49646 42702 49698 42754
rect 50094 42702 50146 42754
rect 50766 42702 50818 42754
rect 50878 42702 50930 42754
rect 55582 42702 55634 42754
rect 17166 42590 17218 42642
rect 20526 42590 20578 42642
rect 23662 42590 23714 42642
rect 24222 42590 24274 42642
rect 29150 42590 29202 42642
rect 30382 42590 30434 42642
rect 31390 42590 31442 42642
rect 35646 42590 35698 42642
rect 35982 42590 36034 42642
rect 41358 42590 41410 42642
rect 42702 42590 42754 42642
rect 43038 42590 43090 42642
rect 46734 42590 46786 42642
rect 50430 42590 50482 42642
rect 19742 42478 19794 42530
rect 20638 42478 20690 42530
rect 20862 42478 20914 42530
rect 23774 42478 23826 42530
rect 23998 42478 24050 42530
rect 24446 42478 24498 42530
rect 25230 42478 25282 42530
rect 27470 42478 27522 42530
rect 28590 42478 28642 42530
rect 30830 42478 30882 42530
rect 30942 42478 30994 42530
rect 31614 42478 31666 42530
rect 32174 42478 32226 42530
rect 33742 42478 33794 42530
rect 36094 42478 36146 42530
rect 39230 42478 39282 42530
rect 43262 42478 43314 42530
rect 43486 42478 43538 42530
rect 45614 42478 45666 42530
rect 45838 42478 45890 42530
rect 46510 42478 46562 42530
rect 46846 42478 46898 42530
rect 50654 42478 50706 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 15598 42142 15650 42194
rect 18286 42142 18338 42194
rect 18846 42142 18898 42194
rect 21646 42142 21698 42194
rect 26126 42142 26178 42194
rect 26350 42142 26402 42194
rect 27918 42142 27970 42194
rect 31502 42142 31554 42194
rect 35198 42142 35250 42194
rect 35870 42142 35922 42194
rect 38670 42142 38722 42194
rect 41470 42142 41522 42194
rect 46286 42142 46338 42194
rect 47182 42142 47234 42194
rect 51774 42142 51826 42194
rect 12014 42030 12066 42082
rect 14254 42030 14306 42082
rect 15822 42030 15874 42082
rect 16830 42030 16882 42082
rect 18734 42030 18786 42082
rect 22878 42030 22930 42082
rect 27358 42030 27410 42082
rect 29262 42030 29314 42082
rect 31726 42030 31778 42082
rect 34190 42030 34242 42082
rect 34414 42030 34466 42082
rect 34638 42030 34690 42082
rect 9662 41918 9714 41970
rect 11566 41918 11618 41970
rect 13246 41918 13298 41970
rect 13918 41918 13970 41970
rect 16046 41918 16098 41970
rect 16606 41918 16658 41970
rect 21982 41918 22034 41970
rect 22654 41918 22706 41970
rect 24222 41918 24274 41970
rect 24782 41918 24834 41970
rect 26014 41918 26066 41970
rect 26574 41918 26626 41970
rect 27022 41918 27074 41970
rect 28030 41918 28082 41970
rect 28702 41918 28754 41970
rect 30270 41918 30322 41970
rect 32174 41918 32226 41970
rect 34750 41918 34802 41970
rect 34862 41918 34914 41970
rect 35310 41918 35362 41970
rect 35534 41918 35586 41970
rect 36206 41918 36258 41970
rect 39006 41918 39058 41970
rect 39790 41918 39842 41970
rect 43822 41918 43874 41970
rect 45390 41918 45442 41970
rect 45614 41918 45666 41970
rect 50654 41918 50706 41970
rect 51102 41918 51154 41970
rect 51438 41918 51490 41970
rect 9998 41806 10050 41858
rect 14030 41806 14082 41858
rect 14814 41806 14866 41858
rect 15150 41806 15202 41858
rect 16158 41806 16210 41858
rect 18398 41806 18450 41858
rect 19854 41806 19906 41858
rect 19966 41806 20018 41858
rect 15262 41694 15314 41746
rect 18062 41694 18114 41746
rect 18846 41694 18898 41746
rect 20414 41806 20466 41858
rect 20974 41806 21026 41858
rect 21422 41806 21474 41858
rect 23214 41806 23266 41858
rect 25566 41806 25618 41858
rect 26462 41806 26514 41858
rect 33182 41806 33234 41858
rect 33630 41806 33682 41858
rect 39678 41806 39730 41858
rect 43934 41806 43986 41858
rect 46622 41806 46674 41858
rect 50206 41806 50258 41858
rect 21310 41694 21362 41746
rect 24558 41694 24610 41746
rect 39902 41694 39954 41746
rect 44494 41694 44546 41746
rect 45838 41694 45890 41746
rect 46846 41694 46898 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 14926 41358 14978 41410
rect 18846 41358 18898 41410
rect 19182 41358 19234 41410
rect 36206 41358 36258 41410
rect 45390 41358 45442 41410
rect 1710 41246 1762 41298
rect 8878 41246 8930 41298
rect 9886 41246 9938 41298
rect 10222 41246 10274 41298
rect 11342 41246 11394 41298
rect 15262 41246 15314 41298
rect 16270 41246 16322 41298
rect 18286 41246 18338 41298
rect 21534 41246 21586 41298
rect 22094 41246 22146 41298
rect 24894 41246 24946 41298
rect 27470 41246 27522 41298
rect 29374 41246 29426 41298
rect 30382 41246 30434 41298
rect 32398 41246 32450 41298
rect 34302 41246 34354 41298
rect 35758 41246 35810 41298
rect 39118 41246 39170 41298
rect 44830 41246 44882 41298
rect 45950 41246 46002 41298
rect 49534 41246 49586 41298
rect 57934 41246 57986 41298
rect 10782 41134 10834 41186
rect 11790 41134 11842 41186
rect 12350 41134 12402 41186
rect 13470 41134 13522 41186
rect 14590 41134 14642 41186
rect 16830 41134 16882 41186
rect 18622 41134 18674 41186
rect 22430 41134 22482 41186
rect 24670 41134 24722 41186
rect 25006 41134 25058 41186
rect 26014 41134 26066 41186
rect 27022 41134 27074 41186
rect 28030 41134 28082 41186
rect 28478 41134 28530 41186
rect 31054 41134 31106 41186
rect 32174 41134 32226 41186
rect 32510 41134 32562 41186
rect 33518 41134 33570 41186
rect 34078 41134 34130 41186
rect 35870 41134 35922 41186
rect 45054 41134 45106 41186
rect 47406 41134 47458 41186
rect 48414 41134 48466 41186
rect 49198 41134 49250 41186
rect 55582 41134 55634 41186
rect 8990 41022 9042 41074
rect 12686 41022 12738 41074
rect 13582 41022 13634 41074
rect 19518 41022 19570 41074
rect 19742 41022 19794 41074
rect 22318 41022 22370 41074
rect 30494 41022 30546 41074
rect 30830 41022 30882 41074
rect 31502 41022 31554 41074
rect 33070 41022 33122 41074
rect 34414 41022 34466 41074
rect 35086 41022 35138 41074
rect 35534 41022 35586 41074
rect 36318 41022 36370 41074
rect 46398 41022 46450 41074
rect 48078 41022 48130 41074
rect 49870 41022 49922 41074
rect 8766 40910 8818 40962
rect 9326 40910 9378 40962
rect 12014 40910 12066 40962
rect 14478 40910 14530 40962
rect 15038 40910 15090 40962
rect 19630 40910 19682 40962
rect 20302 40910 20354 40962
rect 20750 40910 20802 40962
rect 29822 40910 29874 40962
rect 30270 40910 30322 40962
rect 39566 40910 39618 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 15262 40574 15314 40626
rect 15486 40574 15538 40626
rect 15710 40574 15762 40626
rect 16718 40574 16770 40626
rect 26238 40574 26290 40626
rect 27246 40574 27298 40626
rect 10670 40462 10722 40514
rect 11118 40462 11170 40514
rect 13246 40462 13298 40514
rect 14814 40462 14866 40514
rect 16270 40462 16322 40514
rect 16494 40462 16546 40514
rect 20078 40518 20130 40570
rect 27470 40574 27522 40626
rect 35646 40574 35698 40626
rect 43486 40574 43538 40626
rect 50430 40574 50482 40626
rect 17726 40462 17778 40514
rect 18062 40462 18114 40514
rect 18286 40462 18338 40514
rect 18734 40462 18786 40514
rect 21534 40462 21586 40514
rect 25342 40462 25394 40514
rect 26798 40462 26850 40514
rect 34302 40462 34354 40514
rect 36542 40462 36594 40514
rect 39006 40462 39058 40514
rect 39454 40462 39506 40514
rect 41246 40462 41298 40514
rect 10222 40350 10274 40402
rect 11006 40350 11058 40402
rect 13358 40350 13410 40402
rect 13694 40350 13746 40402
rect 14254 40350 14306 40402
rect 16830 40350 16882 40402
rect 19182 40350 19234 40402
rect 19854 40350 19906 40402
rect 20302 40350 20354 40402
rect 20638 40350 20690 40402
rect 21198 40350 21250 40402
rect 24110 40350 24162 40402
rect 24670 40350 24722 40402
rect 25230 40350 25282 40402
rect 26126 40350 26178 40402
rect 27582 40350 27634 40402
rect 27918 40350 27970 40402
rect 28702 40350 28754 40402
rect 29822 40350 29874 40402
rect 30942 40350 30994 40402
rect 32286 40350 32338 40402
rect 33294 40350 33346 40402
rect 37774 40350 37826 40402
rect 39118 40350 39170 40402
rect 41582 40350 41634 40402
rect 42478 40350 42530 40402
rect 44046 40350 44098 40402
rect 49086 40350 49138 40402
rect 49534 40350 49586 40402
rect 49758 40350 49810 40402
rect 50094 40350 50146 40402
rect 14702 40238 14754 40290
rect 15598 40238 15650 40290
rect 17390 40238 17442 40290
rect 17502 40238 17554 40290
rect 18398 40238 18450 40290
rect 18958 40238 19010 40290
rect 20190 40238 20242 40290
rect 22430 40238 22482 40290
rect 26686 40238 26738 40290
rect 27022 40238 27074 40290
rect 35086 40238 35138 40290
rect 36318 40238 36370 40290
rect 38446 40238 38498 40290
rect 43150 40238 43202 40290
rect 31838 40126 31890 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 16830 39790 16882 39842
rect 34190 39790 34242 39842
rect 37550 39790 37602 39842
rect 45726 39790 45778 39842
rect 9102 39678 9154 39730
rect 9886 39678 9938 39730
rect 11342 39678 11394 39730
rect 12798 39678 12850 39730
rect 13582 39678 13634 39730
rect 14478 39678 14530 39730
rect 19406 39678 19458 39730
rect 19966 39678 20018 39730
rect 22766 39678 22818 39730
rect 24110 39678 24162 39730
rect 25342 39678 25394 39730
rect 28478 39678 28530 39730
rect 30830 39678 30882 39730
rect 38222 39678 38274 39730
rect 39566 39678 39618 39730
rect 8542 39566 8594 39618
rect 9438 39566 9490 39618
rect 11790 39566 11842 39618
rect 12686 39566 12738 39618
rect 12910 39566 12962 39618
rect 15150 39566 15202 39618
rect 16382 39566 16434 39618
rect 17278 39566 17330 39618
rect 18062 39566 18114 39618
rect 19182 39566 19234 39618
rect 20190 39566 20242 39618
rect 20526 39566 20578 39618
rect 21646 39566 21698 39618
rect 23886 39566 23938 39618
rect 24222 39566 24274 39618
rect 25566 39566 25618 39618
rect 25790 39566 25842 39618
rect 26350 39566 26402 39618
rect 27358 39566 27410 39618
rect 27582 39566 27634 39618
rect 28366 39566 28418 39618
rect 29262 39566 29314 39618
rect 29598 39566 29650 39618
rect 30382 39566 30434 39618
rect 31166 39566 31218 39618
rect 31390 39566 31442 39618
rect 32958 39566 33010 39618
rect 33182 39566 33234 39618
rect 35982 39566 36034 39618
rect 36318 39566 36370 39618
rect 37214 39566 37266 39618
rect 38558 39566 38610 39618
rect 39118 39566 39170 39618
rect 40574 39566 40626 39618
rect 41134 39566 41186 39618
rect 41582 39566 41634 39618
rect 42142 39566 42194 39618
rect 42366 39566 42418 39618
rect 43150 39566 43202 39618
rect 43374 39566 43426 39618
rect 43486 39566 43538 39618
rect 43934 39566 43986 39618
rect 45390 39566 45442 39618
rect 46398 39566 46450 39618
rect 46622 39566 46674 39618
rect 46846 39566 46898 39618
rect 12014 39454 12066 39506
rect 17838 39454 17890 39506
rect 18958 39454 19010 39506
rect 19518 39454 19570 39506
rect 20750 39454 20802 39506
rect 21310 39454 21362 39506
rect 21422 39454 21474 39506
rect 24894 39454 24946 39506
rect 25230 39454 25282 39506
rect 26126 39454 26178 39506
rect 29374 39454 29426 39506
rect 36430 39454 36482 39506
rect 37438 39454 37490 39506
rect 39230 39454 39282 39506
rect 40238 39454 40290 39506
rect 42702 39454 42754 39506
rect 45166 39454 45218 39506
rect 10782 39342 10834 39394
rect 12462 39342 12514 39394
rect 14030 39342 14082 39394
rect 20862 39342 20914 39394
rect 23214 39342 23266 39394
rect 26910 39342 26962 39394
rect 29822 39342 29874 39394
rect 41022 39342 41074 39394
rect 41470 39342 41522 39394
rect 41694 39342 41746 39394
rect 46510 39342 46562 39394
rect 58158 39342 58210 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 8654 39006 8706 39058
rect 11454 39006 11506 39058
rect 14590 39006 14642 39058
rect 17390 39006 17442 39058
rect 17726 39006 17778 39058
rect 22766 39006 22818 39058
rect 29598 39006 29650 39058
rect 31166 39006 31218 39058
rect 31278 39006 31330 39058
rect 33294 39006 33346 39058
rect 34414 39006 34466 39058
rect 39790 39006 39842 39058
rect 41246 39006 41298 39058
rect 41694 39006 41746 39058
rect 42142 39006 42194 39058
rect 46286 39006 46338 39058
rect 10894 38894 10946 38946
rect 12126 38894 12178 38946
rect 15150 38894 15202 38946
rect 16718 38894 16770 38946
rect 20862 38894 20914 38946
rect 24110 38894 24162 38946
rect 29150 38894 29202 38946
rect 30046 38894 30098 38946
rect 33518 38894 33570 38946
rect 42254 38894 42306 38946
rect 43038 38894 43090 38946
rect 47518 38894 47570 38946
rect 58158 38894 58210 38946
rect 10446 38782 10498 38834
rect 11902 38782 11954 38834
rect 13470 38782 13522 38834
rect 15710 38782 15762 38834
rect 16158 38782 16210 38834
rect 19966 38782 20018 38834
rect 20414 38782 20466 38834
rect 21422 38782 21474 38834
rect 22990 38782 23042 38834
rect 23438 38782 23490 38834
rect 23662 38782 23714 38834
rect 23998 38782 24050 38834
rect 26350 38782 26402 38834
rect 27806 38782 27858 38834
rect 28142 38782 28194 38834
rect 30606 38782 30658 38834
rect 31054 38782 31106 38834
rect 31614 38782 31666 38834
rect 34638 38782 34690 38834
rect 43150 38782 43202 38834
rect 43486 38782 43538 38834
rect 45838 38782 45890 38834
rect 46398 38782 46450 38834
rect 46510 38782 46562 38834
rect 46846 38782 46898 38834
rect 47406 38782 47458 38834
rect 8766 38670 8818 38722
rect 13246 38670 13298 38722
rect 16046 38670 16098 38722
rect 21534 38670 21586 38722
rect 23214 38670 23266 38722
rect 24670 38670 24722 38722
rect 25342 38670 25394 38722
rect 30270 38670 30322 38722
rect 33406 38670 33458 38722
rect 41582 38670 41634 38722
rect 43262 38670 43314 38722
rect 47854 38670 47906 38722
rect 34302 38558 34354 38610
rect 42142 38558 42194 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 15934 38222 15986 38274
rect 23886 38222 23938 38274
rect 29710 38222 29762 38274
rect 37550 38222 37602 38274
rect 37774 38222 37826 38274
rect 12910 38110 12962 38162
rect 21646 38110 21698 38162
rect 22878 38110 22930 38162
rect 25006 38110 25058 38162
rect 26014 38110 26066 38162
rect 28254 38110 28306 38162
rect 31166 38110 31218 38162
rect 32286 38110 32338 38162
rect 46846 38110 46898 38162
rect 57934 38110 57986 38162
rect 9662 37998 9714 38050
rect 11006 37998 11058 38050
rect 12350 37998 12402 38050
rect 13806 37998 13858 38050
rect 14030 37998 14082 38050
rect 14478 37998 14530 38050
rect 16494 37998 16546 38050
rect 17166 37998 17218 38050
rect 19294 37998 19346 38050
rect 19518 37998 19570 38050
rect 24110 37998 24162 38050
rect 24894 37998 24946 38050
rect 25118 37998 25170 38050
rect 25342 37998 25394 38050
rect 26126 37998 26178 38050
rect 27918 37998 27970 38050
rect 29598 37998 29650 38050
rect 31614 37998 31666 38050
rect 32622 37998 32674 38050
rect 32846 37998 32898 38050
rect 33182 37998 33234 38050
rect 33406 37998 33458 38050
rect 33966 37998 34018 38050
rect 34526 37998 34578 38050
rect 35086 37998 35138 38050
rect 35198 37998 35250 38050
rect 35422 37998 35474 38050
rect 42814 37998 42866 38050
rect 48190 37998 48242 38050
rect 55582 37998 55634 38050
rect 11118 37886 11170 37938
rect 11454 37886 11506 37938
rect 12126 37886 12178 37938
rect 16606 37886 16658 37938
rect 17390 37886 17442 37938
rect 19630 37886 19682 37938
rect 24334 37886 24386 37938
rect 25566 37886 25618 37938
rect 25902 37886 25954 37938
rect 29262 37886 29314 37938
rect 29710 37886 29762 37938
rect 31950 37886 32002 37938
rect 34638 37886 34690 37938
rect 34974 37886 35026 37938
rect 36990 37886 37042 37938
rect 37886 37886 37938 37938
rect 42478 37886 42530 37938
rect 47182 37886 47234 37938
rect 48862 37886 48914 37938
rect 49198 37886 49250 37938
rect 49534 37886 49586 37938
rect 1710 37774 1762 37826
rect 9102 37774 9154 37826
rect 22206 37774 22258 37826
rect 23214 37774 23266 37826
rect 23550 37774 23602 37826
rect 23774 37774 23826 37826
rect 24446 37774 24498 37826
rect 24670 37774 24722 37826
rect 26350 37774 26402 37826
rect 26798 37774 26850 37826
rect 27470 37774 27522 37826
rect 30718 37774 30770 37826
rect 31726 37774 31778 37826
rect 37214 37774 37266 37826
rect 37438 37774 37490 37826
rect 42590 37774 42642 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 18062 37438 18114 37490
rect 20414 37438 20466 37490
rect 34302 37438 34354 37490
rect 35646 37438 35698 37490
rect 37214 37438 37266 37490
rect 41918 37438 41970 37490
rect 43934 37438 43986 37490
rect 47294 37438 47346 37490
rect 8990 37326 9042 37378
rect 12462 37326 12514 37378
rect 18958 37326 19010 37378
rect 21198 37326 21250 37378
rect 25566 37326 25618 37378
rect 36878 37326 36930 37378
rect 36990 37326 37042 37378
rect 38558 37326 38610 37378
rect 39342 37326 39394 37378
rect 41134 37326 41186 37378
rect 46734 37326 46786 37378
rect 7870 37214 7922 37266
rect 8318 37214 8370 37266
rect 9662 37214 9714 37266
rect 10894 37214 10946 37266
rect 12798 37214 12850 37266
rect 13806 37214 13858 37266
rect 16046 37214 16098 37266
rect 18174 37214 18226 37266
rect 19854 37214 19906 37266
rect 21870 37214 21922 37266
rect 22766 37214 22818 37266
rect 24334 37214 24386 37266
rect 25230 37214 25282 37266
rect 27022 37214 27074 37266
rect 29262 37214 29314 37266
rect 31054 37214 31106 37266
rect 31278 37214 31330 37266
rect 31502 37214 31554 37266
rect 31614 37214 31666 37266
rect 33742 37214 33794 37266
rect 34190 37214 34242 37266
rect 34414 37214 34466 37266
rect 35198 37214 35250 37266
rect 37998 37214 38050 37266
rect 39230 37214 39282 37266
rect 39566 37214 39618 37266
rect 39790 37214 39842 37266
rect 40910 37214 40962 37266
rect 41806 37214 41858 37266
rect 43710 37214 43762 37266
rect 44382 37214 44434 37266
rect 13694 37102 13746 37154
rect 16830 37102 16882 37154
rect 21534 37102 21586 37154
rect 26350 37102 26402 37154
rect 28030 37102 28082 37154
rect 29822 37102 29874 37154
rect 30270 37102 30322 37154
rect 30718 37102 30770 37154
rect 31390 37102 31442 37154
rect 34750 37102 34802 37154
rect 37774 37102 37826 37154
rect 40014 37102 40066 37154
rect 43822 37102 43874 37154
rect 46958 37102 47010 37154
rect 12910 36990 12962 37042
rect 14366 36990 14418 37042
rect 34974 36990 35026 37042
rect 40126 36990 40178 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 17614 36654 17666 36706
rect 25118 36654 25170 36706
rect 28478 36654 28530 36706
rect 44382 36654 44434 36706
rect 47406 36654 47458 36706
rect 11230 36542 11282 36594
rect 12462 36542 12514 36594
rect 13806 36542 13858 36594
rect 18734 36542 18786 36594
rect 18958 36542 19010 36594
rect 20078 36542 20130 36594
rect 26798 36542 26850 36594
rect 29262 36542 29314 36594
rect 30270 36542 30322 36594
rect 34302 36542 34354 36594
rect 39454 36542 39506 36594
rect 45614 36542 45666 36594
rect 47070 36542 47122 36594
rect 57934 36542 57986 36594
rect 11006 36430 11058 36482
rect 14926 36430 14978 36482
rect 15822 36430 15874 36482
rect 16494 36430 16546 36482
rect 16718 36430 16770 36482
rect 17390 36430 17442 36482
rect 18622 36430 18674 36482
rect 19294 36430 19346 36482
rect 20190 36430 20242 36482
rect 21534 36430 21586 36482
rect 22766 36430 22818 36482
rect 23550 36430 23602 36482
rect 24558 36430 24610 36482
rect 26014 36430 26066 36482
rect 27134 36430 27186 36482
rect 27918 36430 27970 36482
rect 28142 36430 28194 36482
rect 29150 36430 29202 36482
rect 30606 36430 30658 36482
rect 31054 36430 31106 36482
rect 32398 36430 32450 36482
rect 32734 36430 32786 36482
rect 33070 36430 33122 36482
rect 35646 36430 35698 36482
rect 37886 36430 37938 36482
rect 39118 36430 39170 36482
rect 40910 36430 40962 36482
rect 42254 36430 42306 36482
rect 42590 36430 42642 36482
rect 42814 36430 42866 36482
rect 44046 36430 44098 36482
rect 45838 36430 45890 36482
rect 46846 36430 46898 36482
rect 55582 36430 55634 36482
rect 9998 36318 10050 36370
rect 14030 36318 14082 36370
rect 19518 36318 19570 36370
rect 20750 36318 20802 36370
rect 29262 36318 29314 36370
rect 34526 36318 34578 36370
rect 37998 36318 38050 36370
rect 38782 36318 38834 36370
rect 39902 36318 39954 36370
rect 41582 36318 41634 36370
rect 41918 36318 41970 36370
rect 42030 36318 42082 36370
rect 43486 36318 43538 36370
rect 43822 36318 43874 36370
rect 46510 36318 46562 36370
rect 9214 36206 9266 36258
rect 11454 36206 11506 36258
rect 12910 36206 12962 36258
rect 44270 36206 44322 36258
rect 44830 36206 44882 36258
rect 45166 36206 45218 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 13246 35870 13298 35922
rect 14590 35870 14642 35922
rect 23550 35870 23602 35922
rect 24222 35870 24274 35922
rect 24446 35870 24498 35922
rect 29038 35870 29090 35922
rect 30606 35870 30658 35922
rect 32174 35870 32226 35922
rect 34190 35870 34242 35922
rect 34862 35870 34914 35922
rect 35534 35870 35586 35922
rect 35646 35870 35698 35922
rect 36878 35870 36930 35922
rect 39678 35870 39730 35922
rect 40014 35870 40066 35922
rect 42702 35870 42754 35922
rect 43038 35870 43090 35922
rect 7870 35758 7922 35810
rect 9550 35758 9602 35810
rect 11342 35758 11394 35810
rect 11678 35758 11730 35810
rect 14142 35758 14194 35810
rect 15710 35758 15762 35810
rect 27582 35758 27634 35810
rect 30158 35758 30210 35810
rect 31726 35758 31778 35810
rect 34526 35758 34578 35810
rect 34638 35758 34690 35810
rect 44494 35758 44546 35810
rect 46734 35758 46786 35810
rect 8766 35646 8818 35698
rect 9998 35646 10050 35698
rect 10782 35646 10834 35698
rect 11902 35646 11954 35698
rect 13694 35646 13746 35698
rect 14590 35646 14642 35698
rect 15262 35646 15314 35698
rect 16046 35646 16098 35698
rect 17726 35646 17778 35698
rect 18510 35646 18562 35698
rect 19406 35646 19458 35698
rect 20974 35646 21026 35698
rect 21422 35646 21474 35698
rect 23214 35646 23266 35698
rect 24670 35646 24722 35698
rect 25342 35646 25394 35698
rect 25566 35646 25618 35698
rect 26686 35646 26738 35698
rect 27470 35646 27522 35698
rect 28926 35646 28978 35698
rect 30942 35646 30994 35698
rect 33854 35646 33906 35698
rect 34974 35646 35026 35698
rect 35422 35646 35474 35698
rect 36206 35646 36258 35698
rect 36430 35646 36482 35698
rect 43598 35646 43650 35698
rect 43934 35646 43986 35698
rect 46510 35646 46562 35698
rect 16606 35534 16658 35586
rect 17502 35534 17554 35586
rect 18062 35534 18114 35586
rect 21870 35534 21922 35586
rect 24558 35534 24610 35586
rect 26238 35534 26290 35586
rect 30606 35534 30658 35586
rect 33630 35534 33682 35586
rect 35982 35534 36034 35586
rect 21758 35422 21810 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 9326 35086 9378 35138
rect 17390 35086 17442 35138
rect 19406 35086 19458 35138
rect 25006 35086 25058 35138
rect 28590 35086 28642 35138
rect 29822 35086 29874 35138
rect 31166 35086 31218 35138
rect 10782 34974 10834 35026
rect 14030 34974 14082 35026
rect 15374 34974 15426 35026
rect 18398 34974 18450 35026
rect 19966 34974 20018 35026
rect 21758 34974 21810 35026
rect 24222 34974 24274 35026
rect 24894 34974 24946 35026
rect 27358 34974 27410 35026
rect 28142 34974 28194 35026
rect 30270 34974 30322 35026
rect 32398 34974 32450 35026
rect 34638 34974 34690 35026
rect 36318 34974 36370 35026
rect 40686 34974 40738 35026
rect 57822 34974 57874 35026
rect 8766 34862 8818 34914
rect 8990 34862 9042 34914
rect 10894 34862 10946 34914
rect 11790 34862 11842 34914
rect 12910 34862 12962 34914
rect 14814 34862 14866 34914
rect 16046 34862 16098 34914
rect 19294 34862 19346 34914
rect 23550 34862 23602 34914
rect 25790 34862 25842 34914
rect 26014 34862 26066 34914
rect 26686 34862 26738 34914
rect 29262 34862 29314 34914
rect 29486 34862 29538 34914
rect 29710 34862 29762 34914
rect 30606 34862 30658 34914
rect 35086 34862 35138 34914
rect 35870 34862 35922 34914
rect 40350 34862 40402 34914
rect 55582 34862 55634 34914
rect 16494 34750 16546 34802
rect 19182 34750 19234 34802
rect 20414 34750 20466 34802
rect 22766 34750 22818 34802
rect 27022 34750 27074 34802
rect 28478 34750 28530 34802
rect 31054 34750 31106 34802
rect 31166 34750 31218 34802
rect 32510 34750 32562 34802
rect 35534 34750 35586 34802
rect 40014 34750 40066 34802
rect 41358 34750 41410 34802
rect 13582 34638 13634 34690
rect 14478 34638 14530 34690
rect 17950 34638 18002 34690
rect 20750 34638 20802 34690
rect 21310 34638 21362 34690
rect 22318 34638 22370 34690
rect 25454 34638 25506 34690
rect 26350 34638 26402 34690
rect 34862 34638 34914 34690
rect 41022 34638 41074 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 14926 34302 14978 34354
rect 15710 34302 15762 34354
rect 16830 34302 16882 34354
rect 17726 34302 17778 34354
rect 19182 34302 19234 34354
rect 33406 34302 33458 34354
rect 33854 34302 33906 34354
rect 38110 34302 38162 34354
rect 41470 34302 41522 34354
rect 43374 34302 43426 34354
rect 44494 34302 44546 34354
rect 10670 34190 10722 34242
rect 14702 34190 14754 34242
rect 19854 34190 19906 34242
rect 24334 34190 24386 34242
rect 24446 34190 24498 34242
rect 24670 34190 24722 34242
rect 31838 34190 31890 34242
rect 33070 34190 33122 34242
rect 37326 34190 37378 34242
rect 58158 34190 58210 34242
rect 4174 34078 4226 34130
rect 8990 34078 9042 34130
rect 9662 34078 9714 34130
rect 10110 34078 10162 34130
rect 11118 34078 11170 34130
rect 12350 34078 12402 34130
rect 13582 34078 13634 34130
rect 14590 34078 14642 34130
rect 16270 34078 16322 34130
rect 18286 34078 18338 34130
rect 18622 34078 18674 34130
rect 18846 34078 18898 34130
rect 20190 34078 20242 34130
rect 22654 34078 22706 34130
rect 23214 34078 23266 34130
rect 26126 34078 26178 34130
rect 28366 34078 28418 34130
rect 28702 34078 28754 34130
rect 29038 34078 29090 34130
rect 30718 34078 30770 34130
rect 32174 34078 32226 34130
rect 34414 34078 34466 34130
rect 34974 34078 35026 34130
rect 39118 34078 39170 34130
rect 39790 34078 39842 34130
rect 40910 34078 40962 34130
rect 41134 34078 41186 34130
rect 43150 34078 43202 34130
rect 43486 34078 43538 34130
rect 44158 34078 44210 34130
rect 44606 34078 44658 34130
rect 4846 33966 4898 34018
rect 8542 33966 8594 34018
rect 11678 33966 11730 34018
rect 15150 33966 15202 34018
rect 20974 33966 21026 34018
rect 25566 33966 25618 34018
rect 26574 33966 26626 34018
rect 31166 33966 31218 34018
rect 39454 33966 39506 34018
rect 1934 33854 1986 33906
rect 15374 33854 15426 33906
rect 23886 33854 23938 33906
rect 24110 33854 24162 33906
rect 30046 33854 30098 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 10446 33518 10498 33570
rect 19518 33518 19570 33570
rect 25678 33518 25730 33570
rect 35198 33518 35250 33570
rect 1934 33406 1986 33458
rect 12238 33406 12290 33458
rect 14814 33406 14866 33458
rect 17838 33406 17890 33458
rect 18062 33406 18114 33458
rect 18622 33406 18674 33458
rect 19294 33406 19346 33458
rect 20302 33406 20354 33458
rect 23214 33406 23266 33458
rect 24670 33406 24722 33458
rect 25342 33406 25394 33458
rect 26238 33406 26290 33458
rect 26798 33406 26850 33458
rect 38110 33518 38162 33570
rect 27134 33406 27186 33458
rect 28142 33406 28194 33458
rect 29822 33406 29874 33458
rect 37438 33406 37490 33458
rect 37774 33406 37826 33458
rect 4286 33294 4338 33346
rect 9998 33294 10050 33346
rect 10558 33294 10610 33346
rect 10782 33294 10834 33346
rect 12686 33294 12738 33346
rect 16606 33294 16658 33346
rect 17054 33294 17106 33346
rect 18510 33294 18562 33346
rect 22094 33294 22146 33346
rect 22654 33294 22706 33346
rect 23438 33294 23490 33346
rect 24222 33294 24274 33346
rect 25454 33294 25506 33346
rect 27582 33294 27634 33346
rect 28478 33294 28530 33346
rect 29374 33294 29426 33346
rect 30382 33294 30434 33346
rect 30942 33294 30994 33346
rect 31502 33294 31554 33346
rect 32174 33294 32226 33346
rect 35646 33294 35698 33346
rect 36990 33294 37042 33346
rect 40014 33294 40066 33346
rect 42142 33294 42194 33346
rect 43038 33294 43090 33346
rect 45054 33294 45106 33346
rect 15598 33182 15650 33234
rect 17278 33182 17330 33234
rect 24558 33182 24610 33234
rect 29150 33182 29202 33234
rect 30718 33182 30770 33234
rect 40350 33182 40402 33234
rect 42926 33182 42978 33234
rect 9438 33070 9490 33122
rect 11230 33070 11282 33122
rect 16494 33070 16546 33122
rect 19294 33070 19346 33122
rect 20750 33070 20802 33122
rect 21758 33070 21810 33122
rect 23662 33070 23714 33122
rect 24782 33070 24834 33122
rect 34414 33070 34466 33122
rect 37998 33070 38050 33122
rect 38782 33070 38834 33122
rect 41918 33070 41970 33122
rect 42702 33070 42754 33122
rect 44830 33070 44882 33122
rect 58158 33070 58210 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 13470 32734 13522 32786
rect 15934 32734 15986 32786
rect 20750 32734 20802 32786
rect 22430 32734 22482 32786
rect 23886 32734 23938 32786
rect 25902 32734 25954 32786
rect 27918 32734 27970 32786
rect 28702 32734 28754 32786
rect 29038 32734 29090 32786
rect 29374 32734 29426 32786
rect 29710 32734 29762 32786
rect 30382 32734 30434 32786
rect 37438 32734 37490 32786
rect 38110 32734 38162 32786
rect 39454 32734 39506 32786
rect 39678 32734 39730 32786
rect 45390 32734 45442 32786
rect 1710 32622 1762 32674
rect 8878 32622 8930 32674
rect 13582 32622 13634 32674
rect 14254 32622 14306 32674
rect 15710 32622 15762 32674
rect 19070 32622 19122 32674
rect 22878 32622 22930 32674
rect 24670 32622 24722 32674
rect 31614 32622 31666 32674
rect 36878 32622 36930 32674
rect 37214 32622 37266 32674
rect 38334 32622 38386 32674
rect 39118 32622 39170 32674
rect 44606 32622 44658 32674
rect 9774 32510 9826 32562
rect 10670 32510 10722 32562
rect 11230 32510 11282 32562
rect 12462 32510 12514 32562
rect 14030 32510 14082 32562
rect 14814 32510 14866 32562
rect 15598 32510 15650 32562
rect 17838 32510 17890 32562
rect 19406 32510 19458 32562
rect 19966 32510 20018 32562
rect 21422 32510 21474 32562
rect 21646 32510 21698 32562
rect 23326 32510 23378 32562
rect 24110 32510 24162 32562
rect 25454 32510 25506 32562
rect 31838 32510 31890 32562
rect 37886 32510 37938 32562
rect 38222 32510 38274 32562
rect 38782 32510 38834 32562
rect 38894 32510 38946 32562
rect 39230 32510 39282 32562
rect 39790 32510 39842 32562
rect 41694 32510 41746 32562
rect 42254 32510 42306 32562
rect 10222 32398 10274 32450
rect 12126 32398 12178 32450
rect 15150 32398 15202 32450
rect 17950 32398 18002 32450
rect 21534 32398 21586 32450
rect 29822 32398 29874 32450
rect 37326 32398 37378 32450
rect 8990 32286 9042 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 24446 31950 24498 32002
rect 40126 31950 40178 32002
rect 1934 31838 1986 31890
rect 10558 31838 10610 31890
rect 11454 31838 11506 31890
rect 14702 31838 14754 31890
rect 18846 31838 18898 31890
rect 21758 31838 21810 31890
rect 22542 31838 22594 31890
rect 23998 31838 24050 31890
rect 29374 31838 29426 31890
rect 4286 31726 4338 31778
rect 9998 31726 10050 31778
rect 10894 31726 10946 31778
rect 11790 31726 11842 31778
rect 14142 31726 14194 31778
rect 12126 31614 12178 31666
rect 21982 31614 22034 31666
rect 23214 31614 23266 31666
rect 24334 31614 24386 31666
rect 25454 31614 25506 31666
rect 38222 31614 38274 31666
rect 4734 31502 4786 31554
rect 22878 31502 22930 31554
rect 24446 31502 24498 31554
rect 25006 31502 25058 31554
rect 25566 31502 25618 31554
rect 25790 31502 25842 31554
rect 26462 31502 26514 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 8542 31166 8594 31218
rect 9102 31166 9154 31218
rect 12350 31166 12402 31218
rect 13358 31166 13410 31218
rect 14478 31166 14530 31218
rect 18286 31166 18338 31218
rect 18958 31166 19010 31218
rect 19742 31166 19794 31218
rect 20302 31166 20354 31218
rect 22206 31166 22258 31218
rect 23438 31166 23490 31218
rect 23550 31166 23602 31218
rect 23774 31166 23826 31218
rect 24446 31166 24498 31218
rect 24670 31166 24722 31218
rect 30158 31166 30210 31218
rect 44606 31166 44658 31218
rect 45278 31166 45330 31218
rect 9550 31054 9602 31106
rect 16718 31054 16770 31106
rect 19630 31054 19682 31106
rect 23886 31054 23938 31106
rect 29374 31054 29426 31106
rect 35870 31054 35922 31106
rect 38894 31054 38946 31106
rect 57822 31054 57874 31106
rect 4286 30942 4338 30994
rect 5630 30942 5682 30994
rect 6078 30942 6130 30994
rect 9774 30942 9826 30994
rect 12574 30942 12626 30994
rect 13022 30942 13074 30994
rect 14814 30942 14866 30994
rect 15822 30942 15874 30994
rect 18062 30942 18114 30994
rect 18174 30942 18226 30994
rect 18734 30942 18786 30994
rect 19182 30942 19234 30994
rect 21310 30942 21362 30994
rect 21758 30942 21810 30994
rect 24222 30942 24274 30994
rect 25790 30942 25842 30994
rect 26574 30942 26626 30994
rect 27022 30942 27074 30994
rect 32958 30942 33010 30994
rect 33518 30942 33570 30994
rect 38670 30942 38722 30994
rect 41694 30942 41746 30994
rect 42254 30942 42306 30994
rect 58158 30942 58210 30994
rect 1934 30830 1986 30882
rect 15710 30830 15762 30882
rect 20974 30830 21026 30882
rect 22318 30830 22370 30882
rect 22766 30830 22818 30882
rect 24670 30830 24722 30882
rect 25342 30830 25394 30882
rect 26238 30830 26290 30882
rect 57598 30830 57650 30882
rect 19742 30718 19794 30770
rect 36654 30718 36706 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 16606 30382 16658 30434
rect 25342 30382 25394 30434
rect 26462 30382 26514 30434
rect 26798 30382 26850 30434
rect 38894 30382 38946 30434
rect 1710 30270 1762 30322
rect 21870 30270 21922 30322
rect 23886 30270 23938 30322
rect 36206 30270 36258 30322
rect 9102 30158 9154 30210
rect 12238 30158 12290 30210
rect 12574 30158 12626 30210
rect 15822 30158 15874 30210
rect 16494 30158 16546 30210
rect 17390 30158 17442 30210
rect 17838 30158 17890 30210
rect 17950 30158 18002 30210
rect 18622 30158 18674 30210
rect 23662 30158 23714 30210
rect 29822 30158 29874 30210
rect 30270 30158 30322 30210
rect 33294 30158 33346 30210
rect 34750 30158 34802 30210
rect 35534 30158 35586 30210
rect 17726 30046 17778 30098
rect 18286 30046 18338 30098
rect 18734 30046 18786 30098
rect 18958 30046 19010 30098
rect 19182 30046 19234 30098
rect 19630 30046 19682 30098
rect 22990 30046 23042 30098
rect 24334 30046 24386 30098
rect 24558 30046 24610 30098
rect 25790 30046 25842 30098
rect 34862 30046 34914 30098
rect 35870 30046 35922 30098
rect 2158 29934 2210 29986
rect 9662 29934 9714 29986
rect 14926 29934 14978 29986
rect 15262 29934 15314 29986
rect 24446 29934 24498 29986
rect 25118 29934 25170 29986
rect 25230 29934 25282 29986
rect 26686 29934 26738 29986
rect 32734 29934 32786 29986
rect 34526 29934 34578 29986
rect 39118 29934 39170 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 11790 29598 11842 29650
rect 19630 29598 19682 29650
rect 23886 29598 23938 29650
rect 24670 29598 24722 29650
rect 25454 29598 25506 29650
rect 28590 29598 28642 29650
rect 29822 29598 29874 29650
rect 38110 29598 38162 29650
rect 39118 29598 39170 29650
rect 39566 29598 39618 29650
rect 33406 29486 33458 29538
rect 44494 29486 44546 29538
rect 4286 29374 4338 29426
rect 12350 29374 12402 29426
rect 22094 29374 22146 29426
rect 22542 29374 22594 29426
rect 24110 29374 24162 29426
rect 28366 29374 28418 29426
rect 30046 29374 30098 29426
rect 33630 29374 33682 29426
rect 34974 29374 35026 29426
rect 35646 29374 35698 29426
rect 38894 29374 38946 29426
rect 41582 29374 41634 29426
rect 42254 29374 42306 29426
rect 12574 29262 12626 29314
rect 13022 29262 13074 29314
rect 18958 29262 19010 29314
rect 27918 29262 27970 29314
rect 39678 29262 39730 29314
rect 1934 29150 1986 29202
rect 19070 29150 19122 29202
rect 23774 29150 23826 29202
rect 38670 29150 38722 29202
rect 45278 29150 45330 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 17054 28814 17106 28866
rect 28478 28814 28530 28866
rect 24446 28702 24498 28754
rect 34302 28702 34354 28754
rect 6302 28590 6354 28642
rect 12686 28590 12738 28642
rect 13470 28590 13522 28642
rect 13918 28590 13970 28642
rect 20414 28590 20466 28642
rect 25006 28590 25058 28642
rect 25342 28590 25394 28642
rect 29150 28590 29202 28642
rect 30046 28590 30098 28642
rect 30382 28590 30434 28642
rect 33518 28590 33570 28642
rect 34078 28590 34130 28642
rect 36990 28590 37042 28642
rect 38558 28590 38610 28642
rect 39006 28590 39058 28642
rect 42590 28590 42642 28642
rect 43934 28590 43986 28642
rect 45054 28590 45106 28642
rect 5966 28478 6018 28530
rect 12910 28478 12962 28530
rect 18398 28478 18450 28530
rect 18510 28478 18562 28530
rect 20638 28478 20690 28530
rect 23550 28478 23602 28530
rect 27694 28478 27746 28530
rect 29486 28478 29538 28530
rect 32734 28478 32786 28530
rect 42926 28478 42978 28530
rect 43150 28478 43202 28530
rect 43374 28478 43426 28530
rect 43486 28478 43538 28530
rect 1710 28366 1762 28418
rect 16382 28366 16434 28418
rect 18734 28366 18786 28418
rect 19182 28366 19234 28418
rect 23214 28366 23266 28418
rect 33742 28366 33794 28418
rect 37326 28366 37378 28418
rect 41582 28366 41634 28418
rect 42142 28366 42194 28418
rect 42814 28366 42866 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2046 28030 2098 28082
rect 9886 28030 9938 28082
rect 23214 28030 23266 28082
rect 24670 28030 24722 28082
rect 25566 28030 25618 28082
rect 26014 28030 26066 28082
rect 27694 28030 27746 28082
rect 31278 28030 31330 28082
rect 35870 28030 35922 28082
rect 36878 28030 36930 28082
rect 38894 28030 38946 28082
rect 44494 28030 44546 28082
rect 8318 27918 8370 27970
rect 17950 27918 18002 27970
rect 18622 27918 18674 27970
rect 22878 27918 22930 27970
rect 26126 27918 26178 27970
rect 29598 27918 29650 27970
rect 46398 27918 46450 27970
rect 54238 27918 54290 27970
rect 1710 27806 1762 27858
rect 5630 27806 5682 27858
rect 6078 27806 6130 27858
rect 9550 27806 9602 27858
rect 18174 27806 18226 27858
rect 18846 27806 18898 27858
rect 19406 27806 19458 27858
rect 25230 27806 25282 27858
rect 27134 27806 27186 27858
rect 28478 27806 28530 27858
rect 30046 27806 30098 27858
rect 30942 27806 30994 27858
rect 33182 27806 33234 27858
rect 33630 27806 33682 27858
rect 36654 27806 36706 27858
rect 37214 27806 37266 27858
rect 38558 27806 38610 27858
rect 39006 27806 39058 27858
rect 39230 27806 39282 27858
rect 41358 27806 41410 27858
rect 42030 27806 42082 27858
rect 47294 27806 47346 27858
rect 49646 27806 49698 27858
rect 50430 27806 50482 27858
rect 50878 27806 50930 27858
rect 51102 27806 51154 27858
rect 51998 27806 52050 27858
rect 52894 27806 52946 27858
rect 53566 27806 53618 27858
rect 53902 27806 53954 27858
rect 2494 27694 2546 27746
rect 24222 27694 24274 27746
rect 26910 27694 26962 27746
rect 28142 27694 28194 27746
rect 30494 27694 30546 27746
rect 31726 27694 31778 27746
rect 45390 27694 45442 27746
rect 45838 27694 45890 27746
rect 47966 27694 48018 27746
rect 49422 27694 49474 27746
rect 49870 27694 49922 27746
rect 50990 27694 51042 27746
rect 51438 27694 51490 27746
rect 53118 27694 53170 27746
rect 9102 27582 9154 27634
rect 18734 27582 18786 27634
rect 19182 27582 19234 27634
rect 26014 27582 26066 27634
rect 27358 27582 27410 27634
rect 45054 27582 45106 27634
rect 50318 27582 50370 27634
rect 51662 27582 51714 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 43262 27246 43314 27298
rect 47406 27246 47458 27298
rect 49086 27246 49138 27298
rect 49758 27246 49810 27298
rect 49982 27246 50034 27298
rect 57934 27246 57986 27298
rect 1934 27134 1986 27186
rect 10334 27134 10386 27186
rect 25678 27134 25730 27186
rect 26686 27134 26738 27186
rect 41022 27134 41074 27186
rect 53118 27134 53170 27186
rect 4286 27022 4338 27074
rect 8878 27022 8930 27074
rect 9662 27022 9714 27074
rect 18398 27022 18450 27074
rect 18734 27022 18786 27074
rect 22766 27022 22818 27074
rect 33294 27022 33346 27074
rect 34078 27022 34130 27074
rect 37998 27022 38050 27074
rect 41470 27022 41522 27074
rect 45614 27022 45666 27074
rect 46846 27022 46898 27074
rect 49086 27022 49138 27074
rect 49534 27022 49586 27074
rect 51774 27022 51826 27074
rect 52558 27022 52610 27074
rect 55582 27022 55634 27074
rect 9214 26910 9266 26962
rect 9886 26910 9938 26962
rect 12462 26910 12514 26962
rect 15038 26910 15090 26962
rect 16046 26910 16098 26962
rect 22654 26910 22706 26962
rect 23326 26910 23378 26962
rect 23438 26910 23490 26962
rect 30830 26910 30882 26962
rect 33518 26910 33570 26962
rect 33854 26910 33906 26962
rect 38222 26910 38274 26962
rect 38894 26910 38946 26962
rect 43486 26910 43538 26962
rect 45838 26910 45890 26962
rect 47070 26910 47122 26962
rect 47294 26910 47346 26962
rect 48750 26910 48802 26962
rect 50094 26910 50146 26962
rect 51438 26910 51490 26962
rect 51662 26910 51714 26962
rect 12126 26798 12178 26850
rect 15262 26798 15314 26850
rect 22878 26798 22930 26850
rect 23662 26798 23714 26850
rect 40686 26798 40738 26850
rect 43374 26798 43426 26850
rect 46174 26798 46226 26850
rect 46286 26798 46338 26850
rect 46398 26798 46450 26850
rect 53006 26798 53058 26850
rect 53230 26798 53282 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 2046 26462 2098 26514
rect 2718 26462 2770 26514
rect 5070 26462 5122 26514
rect 36542 26462 36594 26514
rect 38558 26462 38610 26514
rect 38782 26462 38834 26514
rect 39566 26462 39618 26514
rect 40238 26462 40290 26514
rect 42142 26462 42194 26514
rect 43374 26462 43426 26514
rect 46510 26462 46562 26514
rect 47070 26462 47122 26514
rect 1710 26350 1762 26402
rect 8206 26350 8258 26402
rect 9662 26350 9714 26402
rect 9998 26350 10050 26402
rect 21198 26350 21250 26402
rect 22542 26350 22594 26402
rect 28366 26350 28418 26402
rect 36206 26350 36258 26402
rect 36878 26350 36930 26402
rect 39678 26350 39730 26402
rect 40350 26350 40402 26402
rect 43038 26350 43090 26402
rect 43150 26350 43202 26402
rect 45838 26350 45890 26402
rect 45950 26350 46002 26402
rect 46286 26350 46338 26402
rect 46622 26350 46674 26402
rect 49758 26350 49810 26402
rect 50318 26350 50370 26402
rect 55022 26350 55074 26402
rect 2382 26238 2434 26290
rect 4398 26238 4450 26290
rect 4846 26238 4898 26290
rect 5518 26238 5570 26290
rect 5966 26238 6018 26290
rect 10446 26238 10498 26290
rect 11230 26238 11282 26290
rect 11790 26238 11842 26290
rect 14030 26238 14082 26290
rect 20078 26238 20130 26290
rect 21646 26238 21698 26290
rect 22990 26238 23042 26290
rect 23774 26238 23826 26290
rect 24222 26238 24274 26290
rect 24334 26238 24386 26290
rect 25902 26238 25954 26290
rect 26126 26238 26178 26290
rect 28254 26238 28306 26290
rect 39230 26238 39282 26290
rect 40014 26238 40066 26290
rect 43710 26238 43762 26290
rect 48862 26238 48914 26290
rect 49086 26238 49138 26290
rect 50206 26238 50258 26290
rect 50542 26238 50594 26290
rect 50766 26238 50818 26290
rect 50990 26238 51042 26290
rect 51998 26238 52050 26290
rect 52334 26238 52386 26290
rect 53006 26238 53058 26290
rect 53678 26238 53730 26290
rect 54350 26238 54402 26290
rect 54686 26238 54738 26290
rect 3166 26126 3218 26178
rect 10782 26126 10834 26178
rect 19630 26126 19682 26178
rect 20414 26126 20466 26178
rect 22094 26126 22146 26178
rect 23326 26126 23378 26178
rect 23998 26126 24050 26178
rect 26014 26126 26066 26178
rect 26910 26126 26962 26178
rect 27470 26126 27522 26178
rect 29038 26126 29090 26178
rect 31054 26126 31106 26178
rect 38222 26126 38274 26178
rect 38670 26126 38722 26178
rect 42702 26126 42754 26178
rect 46958 26126 47010 26178
rect 53566 26126 53618 26178
rect 8990 26014 9042 26066
rect 15038 26014 15090 26066
rect 25342 26014 25394 26066
rect 28366 26014 28418 26066
rect 36990 26014 37042 26066
rect 39454 26014 39506 26066
rect 45950 26014 46002 26066
rect 50766 26014 50818 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 22542 25678 22594 25730
rect 22878 25678 22930 25730
rect 29710 25678 29762 25730
rect 52782 25678 52834 25730
rect 57934 25678 57986 25730
rect 2494 25566 2546 25618
rect 5742 25566 5794 25618
rect 15262 25566 15314 25618
rect 20302 25566 20354 25618
rect 20414 25566 20466 25618
rect 21422 25566 21474 25618
rect 23102 25566 23154 25618
rect 23774 25566 23826 25618
rect 24670 25566 24722 25618
rect 30830 25566 30882 25618
rect 35534 25566 35586 25618
rect 37886 25566 37938 25618
rect 42590 25566 42642 25618
rect 43486 25566 43538 25618
rect 47182 25566 47234 25618
rect 51550 25566 51602 25618
rect 52670 25566 52722 25618
rect 4174 25454 4226 25506
rect 5070 25454 5122 25506
rect 6526 25454 6578 25506
rect 8766 25454 8818 25506
rect 9214 25454 9266 25506
rect 11342 25454 11394 25506
rect 14030 25454 14082 25506
rect 14478 25454 14530 25506
rect 17838 25454 17890 25506
rect 18286 25454 18338 25506
rect 18734 25454 18786 25506
rect 20638 25454 20690 25506
rect 25342 25454 25394 25506
rect 27918 25454 27970 25506
rect 29486 25454 29538 25506
rect 29934 25454 29986 25506
rect 30382 25454 30434 25506
rect 31278 25454 31330 25506
rect 31502 25454 31554 25506
rect 32846 25454 32898 25506
rect 33406 25454 33458 25506
rect 33742 25454 33794 25506
rect 34078 25454 34130 25506
rect 35198 25454 35250 25506
rect 39006 25454 39058 25506
rect 39566 25454 39618 25506
rect 42366 25454 42418 25506
rect 42702 25454 42754 25506
rect 43038 25454 43090 25506
rect 46286 25454 46338 25506
rect 46510 25454 46562 25506
rect 50654 25454 50706 25506
rect 50878 25454 50930 25506
rect 55582 25454 55634 25506
rect 1710 25342 1762 25394
rect 2046 25342 2098 25394
rect 4398 25342 4450 25394
rect 6190 25342 6242 25394
rect 15374 25342 15426 25394
rect 16046 25342 16098 25394
rect 16606 25342 16658 25394
rect 24782 25342 24834 25394
rect 27582 25342 27634 25394
rect 28254 25342 28306 25394
rect 32062 25342 32114 25394
rect 40238 25342 40290 25394
rect 43374 25342 43426 25394
rect 2942 25230 2994 25282
rect 4734 25230 4786 25282
rect 12462 25230 12514 25282
rect 17614 25230 17666 25282
rect 19406 25230 19458 25282
rect 25006 25230 25058 25282
rect 27246 25230 27298 25282
rect 27694 25230 27746 25282
rect 28590 25230 28642 25282
rect 29038 25230 29090 25282
rect 34302 25230 34354 25282
rect 34638 25230 34690 25282
rect 37326 25230 37378 25282
rect 43598 25230 43650 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 20862 24894 20914 24946
rect 25790 24894 25842 24946
rect 34190 24894 34242 24946
rect 42142 24894 42194 24946
rect 48862 24894 48914 24946
rect 53006 24894 53058 24946
rect 19294 24782 19346 24834
rect 23662 24782 23714 24834
rect 4286 24670 4338 24722
rect 5070 24670 5122 24722
rect 5518 24670 5570 24722
rect 7758 24670 7810 24722
rect 14142 24670 14194 24722
rect 15262 24670 15314 24722
rect 16382 24670 16434 24722
rect 17390 24670 17442 24722
rect 17838 24670 17890 24722
rect 12686 24558 12738 24610
rect 13918 24558 13970 24610
rect 18510 24558 18562 24610
rect 19070 24558 19122 24610
rect 1934 24446 1986 24498
rect 8766 24446 8818 24498
rect 16270 24446 16322 24498
rect 18734 24446 18786 24498
rect 29822 24782 29874 24834
rect 33630 24782 33682 24834
rect 34414 24782 34466 24834
rect 35646 24782 35698 24834
rect 41806 24782 41858 24834
rect 43374 24782 43426 24834
rect 49646 24782 49698 24834
rect 19854 24670 19906 24722
rect 23102 24670 23154 24722
rect 26014 24670 26066 24722
rect 26910 24670 26962 24722
rect 28142 24670 28194 24722
rect 28478 24670 28530 24722
rect 30718 24670 30770 24722
rect 30830 24670 30882 24722
rect 31166 24670 31218 24722
rect 32062 24670 32114 24722
rect 33294 24670 33346 24722
rect 33854 24670 33906 24722
rect 35086 24670 35138 24722
rect 35422 24670 35474 24722
rect 43150 24670 43202 24722
rect 44718 24670 44770 24722
rect 46286 24670 46338 24722
rect 47070 24670 47122 24722
rect 48750 24670 48802 24722
rect 48974 24670 49026 24722
rect 49422 24670 49474 24722
rect 52894 24670 52946 24722
rect 53230 24670 53282 24722
rect 53902 24670 53954 24722
rect 19518 24558 19570 24610
rect 20414 24558 20466 24610
rect 22878 24558 22930 24610
rect 25342 24558 25394 24610
rect 25678 24558 25730 24610
rect 26462 24558 26514 24610
rect 28702 24558 28754 24610
rect 31054 24558 31106 24610
rect 31726 24558 31778 24610
rect 34526 24558 34578 24610
rect 34862 24558 34914 24610
rect 36430 24558 36482 24610
rect 36990 24558 37042 24610
rect 44382 24558 44434 24610
rect 23326 24446 23378 24498
rect 23550 24446 23602 24498
rect 28478 24446 28530 24498
rect 29934 24446 29986 24498
rect 34638 24446 34690 24498
rect 34974 24446 35026 24498
rect 35758 24446 35810 24498
rect 36318 24446 36370 24498
rect 36990 24446 37042 24498
rect 49758 24446 49810 24498
rect 55358 24446 55410 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 18286 24110 18338 24162
rect 19518 24110 19570 24162
rect 35646 24110 35698 24162
rect 43150 24110 43202 24162
rect 43486 24110 43538 24162
rect 46846 24110 46898 24162
rect 53678 24110 53730 24162
rect 57934 24110 57986 24162
rect 1934 23998 1986 24050
rect 9550 23998 9602 24050
rect 10446 23998 10498 24050
rect 10894 23998 10946 24050
rect 11902 23998 11954 24050
rect 15934 23998 15986 24050
rect 16270 23998 16322 24050
rect 25230 23998 25282 24050
rect 28366 23998 28418 24050
rect 30046 23998 30098 24050
rect 32958 23998 33010 24050
rect 42478 23998 42530 24050
rect 45614 23998 45666 24050
rect 46958 23998 47010 24050
rect 48190 23998 48242 24050
rect 49310 23998 49362 24050
rect 53342 23998 53394 24050
rect 4286 23886 4338 23938
rect 5966 23886 6018 23938
rect 11230 23886 11282 23938
rect 13918 23886 13970 23938
rect 14366 23886 14418 23938
rect 14926 23886 14978 23938
rect 15374 23886 15426 23938
rect 16494 23886 16546 23938
rect 18622 23886 18674 23938
rect 19294 23886 19346 23938
rect 22990 23886 23042 23938
rect 23550 23886 23602 23938
rect 26126 23886 26178 23938
rect 27134 23886 27186 23938
rect 28142 23886 28194 23938
rect 30494 23886 30546 23938
rect 30942 23886 30994 23938
rect 31726 23886 31778 23938
rect 33406 23886 33458 23938
rect 34750 23886 34802 23938
rect 35758 23886 35810 23938
rect 36206 23886 36258 23938
rect 37102 23886 37154 23938
rect 38782 23886 38834 23938
rect 40798 23886 40850 23938
rect 45166 23886 45218 23938
rect 46062 23886 46114 23938
rect 46734 23886 46786 23938
rect 47966 23886 48018 23938
rect 48862 23886 48914 23938
rect 49758 23886 49810 23938
rect 52894 23886 52946 23938
rect 53454 23886 53506 23938
rect 54686 23886 54738 23938
rect 55582 23886 55634 23938
rect 5630 23774 5682 23826
rect 22878 23774 22930 23826
rect 23774 23774 23826 23826
rect 25006 23774 25058 23826
rect 25566 23774 25618 23826
rect 27582 23774 27634 23826
rect 28030 23774 28082 23826
rect 30270 23774 30322 23826
rect 31838 23774 31890 23826
rect 37886 23774 37938 23826
rect 40350 23774 40402 23826
rect 44830 23774 44882 23826
rect 50206 23774 50258 23826
rect 54462 23774 54514 23826
rect 9102 23662 9154 23714
rect 12350 23662 12402 23714
rect 12798 23662 12850 23714
rect 15038 23662 15090 23714
rect 19854 23662 19906 23714
rect 20526 23662 20578 23714
rect 21534 23662 21586 23714
rect 21982 23662 22034 23714
rect 22654 23662 22706 23714
rect 23102 23662 23154 23714
rect 24334 23662 24386 23714
rect 25342 23662 25394 23714
rect 29486 23662 29538 23714
rect 30606 23662 30658 23714
rect 30718 23662 30770 23714
rect 35646 23662 35698 23714
rect 41246 23662 41298 23714
rect 42030 23662 42082 23714
rect 42590 23662 42642 23714
rect 43374 23662 43426 23714
rect 44270 23662 44322 23714
rect 44942 23662 44994 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 12462 23326 12514 23378
rect 17390 23326 17442 23378
rect 18510 23326 18562 23378
rect 20974 23326 21026 23378
rect 21422 23326 21474 23378
rect 24558 23326 24610 23378
rect 26910 23326 26962 23378
rect 34414 23326 34466 23378
rect 35422 23326 35474 23378
rect 36206 23326 36258 23378
rect 36766 23326 36818 23378
rect 36878 23326 36930 23378
rect 38558 23326 38610 23378
rect 44382 23326 44434 23378
rect 49534 23326 49586 23378
rect 51438 23326 51490 23378
rect 52222 23326 52274 23378
rect 52670 23326 52722 23378
rect 53006 23326 53058 23378
rect 8990 23214 9042 23266
rect 12014 23214 12066 23266
rect 12574 23214 12626 23266
rect 13694 23214 13746 23266
rect 25566 23214 25618 23266
rect 32510 23214 32562 23266
rect 37662 23214 37714 23266
rect 37998 23214 38050 23266
rect 41022 23214 41074 23266
rect 41806 23214 41858 23266
rect 42366 23214 42418 23266
rect 44830 23214 44882 23266
rect 49198 23214 49250 23266
rect 49310 23214 49362 23266
rect 51102 23214 51154 23266
rect 51214 23214 51266 23266
rect 51662 23214 51714 23266
rect 54462 23214 54514 23266
rect 4286 23102 4338 23154
rect 7870 23102 7922 23154
rect 8318 23102 8370 23154
rect 8766 23102 8818 23154
rect 10110 23102 10162 23154
rect 10558 23102 10610 23154
rect 11454 23102 11506 23154
rect 13358 23102 13410 23154
rect 16270 23102 16322 23154
rect 16718 23102 16770 23154
rect 19854 23102 19906 23154
rect 20302 23102 20354 23154
rect 20638 23102 20690 23154
rect 22766 23102 22818 23154
rect 26350 23102 26402 23154
rect 26686 23102 26738 23154
rect 27022 23102 27074 23154
rect 27470 23102 27522 23154
rect 27694 23102 27746 23154
rect 28366 23102 28418 23154
rect 28590 23102 28642 23154
rect 29598 23102 29650 23154
rect 29934 23102 29986 23154
rect 30382 23102 30434 23154
rect 30942 23102 30994 23154
rect 31390 23102 31442 23154
rect 31502 23102 31554 23154
rect 31614 23102 31666 23154
rect 34190 23102 34242 23154
rect 34302 23102 34354 23154
rect 34526 23102 34578 23154
rect 34750 23102 34802 23154
rect 40126 23102 40178 23154
rect 40910 23102 40962 23154
rect 42702 23102 42754 23154
rect 44046 23102 44098 23154
rect 44158 23102 44210 23154
rect 44494 23102 44546 23154
rect 45390 23102 45442 23154
rect 51886 23102 51938 23154
rect 52894 23102 52946 23154
rect 53118 23102 53170 23154
rect 53790 23102 53842 23154
rect 7982 22990 8034 23042
rect 9774 22990 9826 23042
rect 11006 22990 11058 23042
rect 14590 22990 14642 23042
rect 17950 22990 18002 23042
rect 19070 22990 19122 23042
rect 19518 22990 19570 23042
rect 21982 22990 22034 23042
rect 22430 22990 22482 23042
rect 1934 22878 1986 22930
rect 11678 22878 11730 22930
rect 21870 22878 21922 22930
rect 22766 22990 22818 23042
rect 23886 22990 23938 23042
rect 25678 22990 25730 23042
rect 26126 22990 26178 23042
rect 32174 22990 32226 23042
rect 33742 22990 33794 23042
rect 39006 22990 39058 23042
rect 42142 22990 42194 23042
rect 43150 22990 43202 23042
rect 45614 22990 45666 23042
rect 47406 22990 47458 23042
rect 54014 22990 54066 23042
rect 25342 22878 25394 22930
rect 28030 22878 28082 22930
rect 30046 22878 30098 22930
rect 36654 22878 36706 22930
rect 38222 22878 38274 22930
rect 39230 22878 39282 22930
rect 39454 22878 39506 22930
rect 39678 22878 39730 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16494 22542 16546 22594
rect 31278 22542 31330 22594
rect 37774 22542 37826 22594
rect 39230 22542 39282 22594
rect 47966 22542 48018 22594
rect 50766 22542 50818 22594
rect 1934 22430 1986 22482
rect 8878 22430 8930 22482
rect 10894 22430 10946 22482
rect 16046 22430 16098 22482
rect 20078 22430 20130 22482
rect 27806 22430 27858 22482
rect 30046 22430 30098 22482
rect 31054 22430 31106 22482
rect 32622 22430 32674 22482
rect 36430 22430 36482 22482
rect 38110 22430 38162 22482
rect 39006 22430 39058 22482
rect 40014 22430 40066 22482
rect 45390 22430 45442 22482
rect 47294 22430 47346 22482
rect 53790 22430 53842 22482
rect 54350 22430 54402 22482
rect 4174 22318 4226 22370
rect 9326 22318 9378 22370
rect 9662 22318 9714 22370
rect 11230 22318 11282 22370
rect 11342 22318 11394 22370
rect 11566 22318 11618 22370
rect 13806 22318 13858 22370
rect 14254 22318 14306 22370
rect 14590 22318 14642 22370
rect 15374 22318 15426 22370
rect 16382 22318 16434 22370
rect 17166 22318 17218 22370
rect 19294 22318 19346 22370
rect 21646 22318 21698 22370
rect 23662 22318 23714 22370
rect 24782 22318 24834 22370
rect 27470 22318 27522 22370
rect 28254 22318 28306 22370
rect 30270 22318 30322 22370
rect 31390 22318 31442 22370
rect 33070 22318 33122 22370
rect 33966 22318 34018 22370
rect 34974 22318 35026 22370
rect 35310 22318 35362 22370
rect 39454 22318 39506 22370
rect 39790 22318 39842 22370
rect 40126 22318 40178 22370
rect 41358 22318 41410 22370
rect 41582 22318 41634 22370
rect 42030 22318 42082 22370
rect 43710 22318 43762 22370
rect 43822 22318 43874 22370
rect 44718 22318 44770 22370
rect 45502 22318 45554 22370
rect 47518 22318 47570 22370
rect 50206 22318 50258 22370
rect 50430 22318 50482 22370
rect 50654 22318 50706 22370
rect 53902 22318 53954 22370
rect 9774 22206 9826 22258
rect 10222 22206 10274 22258
rect 12126 22206 12178 22258
rect 15150 22206 15202 22258
rect 17278 22206 17330 22258
rect 18174 22206 18226 22258
rect 18286 22206 18338 22258
rect 20526 22206 20578 22258
rect 21982 22206 22034 22258
rect 25454 22206 25506 22258
rect 26126 22206 26178 22258
rect 27134 22206 27186 22258
rect 27806 22206 27858 22258
rect 32846 22206 32898 22258
rect 34302 22206 34354 22258
rect 34526 22206 34578 22258
rect 35534 22206 35586 22258
rect 37998 22206 38050 22258
rect 41806 22206 41858 22258
rect 42142 22206 42194 22258
rect 46174 22206 46226 22258
rect 53566 22206 53618 22258
rect 54238 22206 54290 22258
rect 54462 22206 54514 22258
rect 8430 22094 8482 22146
rect 12910 22094 12962 22146
rect 17502 22094 17554 22146
rect 18510 22094 18562 22146
rect 25230 22094 25282 22146
rect 25790 22094 25842 22146
rect 29374 22094 29426 22146
rect 35422 22094 35474 22146
rect 39902 22094 39954 22146
rect 43038 22094 43090 22146
rect 43374 22094 43426 22146
rect 43934 22094 43986 22146
rect 44158 22094 44210 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 6302 21758 6354 21810
rect 10782 21758 10834 21810
rect 16046 21758 16098 21810
rect 17390 21758 17442 21810
rect 19294 21758 19346 21810
rect 21758 21758 21810 21810
rect 21982 21758 22034 21810
rect 22878 21758 22930 21810
rect 22990 21758 23042 21810
rect 25342 21758 25394 21810
rect 27470 21758 27522 21810
rect 27694 21758 27746 21810
rect 32622 21758 32674 21810
rect 33406 21758 33458 21810
rect 34974 21758 35026 21810
rect 42814 21758 42866 21810
rect 44046 21758 44098 21810
rect 47518 21758 47570 21810
rect 47630 21758 47682 21810
rect 47742 21758 47794 21810
rect 6974 21646 7026 21698
rect 16830 21646 16882 21698
rect 20750 21646 20802 21698
rect 21646 21646 21698 21698
rect 22206 21646 22258 21698
rect 22318 21646 22370 21698
rect 26686 21646 26738 21698
rect 27358 21646 27410 21698
rect 29150 21646 29202 21698
rect 32398 21646 32450 21698
rect 33070 21646 33122 21698
rect 34750 21646 34802 21698
rect 36878 21646 36930 21698
rect 37550 21646 37602 21698
rect 41022 21646 41074 21698
rect 42254 21646 42306 21698
rect 44158 21646 44210 21698
rect 44830 21646 44882 21698
rect 46734 21646 46786 21698
rect 49422 21646 49474 21698
rect 54014 21646 54066 21698
rect 54574 21646 54626 21698
rect 4286 21534 4338 21586
rect 5966 21534 6018 21586
rect 6750 21534 6802 21586
rect 11566 21534 11618 21586
rect 14142 21534 14194 21586
rect 15150 21534 15202 21586
rect 16494 21534 16546 21586
rect 17950 21534 18002 21586
rect 19630 21534 19682 21586
rect 22654 21534 22706 21586
rect 23102 21534 23154 21586
rect 23326 21534 23378 21586
rect 24110 21534 24162 21586
rect 24334 21534 24386 21586
rect 24670 21534 24722 21586
rect 25790 21534 25842 21586
rect 26126 21534 26178 21586
rect 28366 21534 28418 21586
rect 28814 21534 28866 21586
rect 29710 21534 29762 21586
rect 30158 21534 30210 21586
rect 30830 21534 30882 21586
rect 31054 21534 31106 21586
rect 32286 21534 32338 21586
rect 34190 21534 34242 21586
rect 34638 21534 34690 21586
rect 35982 21534 36034 21586
rect 36206 21534 36258 21586
rect 37326 21534 37378 21586
rect 38110 21534 38162 21586
rect 42142 21534 42194 21586
rect 42814 21534 42866 21586
rect 43486 21534 43538 21586
rect 43710 21534 43762 21586
rect 44382 21534 44434 21586
rect 46846 21534 46898 21586
rect 47070 21534 47122 21586
rect 49758 21534 49810 21586
rect 50878 21534 50930 21586
rect 53118 21534 53170 21586
rect 1934 21422 1986 21474
rect 12686 21422 12738 21474
rect 13246 21422 13298 21474
rect 13806 21422 13858 21474
rect 14702 21422 14754 21474
rect 15598 21422 15650 21474
rect 18510 21422 18562 21474
rect 18734 21422 18786 21474
rect 21422 21422 21474 21474
rect 23774 21422 23826 21474
rect 24222 21422 24274 21474
rect 26574 21422 26626 21474
rect 28030 21422 28082 21474
rect 30046 21422 30098 21474
rect 33854 21422 33906 21474
rect 41246 21422 41298 21474
rect 51662 21422 51714 21474
rect 53342 21422 53394 21474
rect 54462 21422 54514 21474
rect 31278 21310 31330 21362
rect 38446 21310 38498 21362
rect 41582 21310 41634 21362
rect 44718 21310 44770 21362
rect 46734 21310 46786 21362
rect 54350 21310 54402 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 30270 20974 30322 21026
rect 37550 20974 37602 21026
rect 47630 20974 47682 21026
rect 49982 20974 50034 21026
rect 11118 20862 11170 20914
rect 12462 20862 12514 20914
rect 22878 20862 22930 20914
rect 23774 20862 23826 20914
rect 27022 20862 27074 20914
rect 31726 20862 31778 20914
rect 36990 20862 37042 20914
rect 38446 20862 38498 20914
rect 39902 20862 39954 20914
rect 47294 20862 47346 20914
rect 49422 20862 49474 20914
rect 50542 20862 50594 20914
rect 51774 20862 51826 20914
rect 57934 20862 57986 20914
rect 5854 20750 5906 20802
rect 7422 20750 7474 20802
rect 7982 20750 8034 20802
rect 12910 20750 12962 20802
rect 14030 20750 14082 20802
rect 15822 20750 15874 20802
rect 17390 20750 17442 20802
rect 19182 20750 19234 20802
rect 20638 20750 20690 20802
rect 24558 20750 24610 20802
rect 25342 20750 25394 20802
rect 27918 20750 27970 20802
rect 31166 20750 31218 20802
rect 31390 20750 31442 20802
rect 33630 20750 33682 20802
rect 35870 20750 35922 20802
rect 37214 20750 37266 20802
rect 37998 20750 38050 20802
rect 41582 20750 41634 20802
rect 42478 20750 42530 20802
rect 46398 20750 46450 20802
rect 46622 20750 46674 20802
rect 49646 20750 49698 20802
rect 50990 20750 51042 20802
rect 51214 20750 51266 20802
rect 54014 20750 54066 20802
rect 54238 20750 54290 20802
rect 55582 20750 55634 20802
rect 11566 20638 11618 20690
rect 14478 20638 14530 20690
rect 15934 20638 15986 20690
rect 17166 20638 17218 20690
rect 19742 20638 19794 20690
rect 20414 20638 20466 20690
rect 20750 20638 20802 20690
rect 21310 20638 21362 20690
rect 21534 20638 21586 20690
rect 21870 20638 21922 20690
rect 22430 20638 22482 20690
rect 24782 20638 24834 20690
rect 25454 20638 25506 20690
rect 25678 20638 25730 20690
rect 30158 20638 30210 20690
rect 31614 20638 31666 20690
rect 33294 20638 33346 20690
rect 35086 20638 35138 20690
rect 36094 20638 36146 20690
rect 40014 20638 40066 20690
rect 40238 20638 40290 20690
rect 40462 20638 40514 20690
rect 40574 20638 40626 20690
rect 41694 20638 41746 20690
rect 45390 20638 45442 20690
rect 47742 20638 47794 20690
rect 50318 20638 50370 20690
rect 54462 20638 54514 20690
rect 54798 20638 54850 20690
rect 55134 20638 55186 20690
rect 6078 20526 6130 20578
rect 6414 20526 6466 20578
rect 6750 20526 6802 20578
rect 7086 20526 7138 20578
rect 7758 20526 7810 20578
rect 10670 20526 10722 20578
rect 12014 20526 12066 20578
rect 13582 20526 13634 20578
rect 18622 20526 18674 20578
rect 21758 20526 21810 20578
rect 22094 20526 22146 20578
rect 22318 20526 22370 20578
rect 23326 20526 23378 20578
rect 26126 20526 26178 20578
rect 26574 20526 26626 20578
rect 27358 20526 27410 20578
rect 28366 20526 28418 20578
rect 29374 20526 29426 20578
rect 29934 20526 29986 20578
rect 30270 20526 30322 20578
rect 31838 20526 31890 20578
rect 32846 20526 32898 20578
rect 39790 20526 39842 20578
rect 42478 20526 42530 20578
rect 44830 20526 44882 20578
rect 50542 20526 50594 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 14478 20190 14530 20242
rect 21086 20190 21138 20242
rect 27582 20190 27634 20242
rect 8094 20078 8146 20130
rect 8654 20078 8706 20130
rect 12350 20078 12402 20130
rect 16830 20078 16882 20130
rect 18398 20078 18450 20130
rect 19070 20078 19122 20130
rect 19518 20078 19570 20130
rect 24334 20078 24386 20130
rect 27134 20078 27186 20130
rect 34078 20078 34130 20130
rect 35870 20078 35922 20130
rect 36542 20078 36594 20130
rect 37438 20078 37490 20130
rect 6414 19966 6466 20018
rect 7086 19966 7138 20018
rect 7310 19966 7362 20018
rect 7982 19966 8034 20018
rect 9998 19966 10050 20018
rect 11342 19966 11394 20018
rect 13134 19966 13186 20018
rect 14590 19966 14642 20018
rect 15486 19966 15538 20018
rect 15710 19966 15762 20018
rect 16382 19966 16434 20018
rect 16606 19966 16658 20018
rect 16942 19966 16994 20018
rect 17726 19966 17778 20018
rect 18734 19966 18786 20018
rect 19742 19966 19794 20018
rect 21198 19966 21250 20018
rect 21534 19966 21586 20018
rect 23326 19966 23378 20018
rect 24110 19966 24162 20018
rect 25342 19966 25394 20018
rect 25678 19966 25730 20018
rect 26238 19966 26290 20018
rect 29038 19966 29090 20018
rect 29262 19966 29314 20018
rect 29710 19966 29762 20018
rect 30382 19966 30434 20018
rect 32398 19966 32450 20018
rect 33518 19966 33570 20018
rect 33742 19966 33794 20018
rect 35198 19966 35250 20018
rect 35646 19966 35698 20018
rect 36318 19966 36370 20018
rect 37998 19966 38050 20018
rect 38222 19966 38274 20018
rect 41582 19966 41634 20018
rect 41918 19966 41970 20018
rect 42142 19966 42194 20018
rect 6078 19854 6130 19906
rect 9662 19854 9714 19906
rect 10446 19854 10498 19906
rect 10558 19854 10610 19906
rect 7646 19742 7698 19794
rect 11006 19854 11058 19906
rect 11902 19854 11954 19906
rect 18062 19854 18114 19906
rect 23774 19854 23826 19906
rect 23998 19854 24050 19906
rect 26798 19854 26850 19906
rect 28142 19854 28194 19906
rect 28478 19854 28530 19906
rect 29150 19854 29202 19906
rect 30046 19854 30098 19906
rect 30942 19854 30994 19906
rect 35422 19854 35474 19906
rect 41806 19854 41858 19906
rect 11118 19742 11170 19794
rect 15150 19742 15202 19794
rect 27358 19742 27410 19794
rect 28478 19742 28530 19794
rect 37102 19742 37154 19794
rect 37886 19742 37938 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14814 19406 14866 19458
rect 19742 19406 19794 19458
rect 21310 19406 21362 19458
rect 21646 19406 21698 19458
rect 24334 19406 24386 19458
rect 30382 19406 30434 19458
rect 34974 19406 35026 19458
rect 41582 19406 41634 19458
rect 41918 19406 41970 19458
rect 17726 19294 17778 19346
rect 20078 19294 20130 19346
rect 21982 19294 22034 19346
rect 27470 19294 27522 19346
rect 28478 19294 28530 19346
rect 30830 19294 30882 19346
rect 31950 19294 32002 19346
rect 35870 19294 35922 19346
rect 46174 19294 46226 19346
rect 47070 19294 47122 19346
rect 51886 19294 51938 19346
rect 5966 19182 6018 19234
rect 6414 19182 6466 19234
rect 8990 19182 9042 19234
rect 9774 19182 9826 19234
rect 10110 19182 10162 19234
rect 10670 19182 10722 19234
rect 11118 19182 11170 19234
rect 13694 19182 13746 19234
rect 15486 19182 15538 19234
rect 17838 19182 17890 19234
rect 18846 19182 18898 19234
rect 19742 19182 19794 19234
rect 22430 19182 22482 19234
rect 24894 19182 24946 19234
rect 25790 19182 25842 19234
rect 26462 19182 26514 19234
rect 26686 19182 26738 19234
rect 26798 19182 26850 19234
rect 27694 19182 27746 19234
rect 29262 19182 29314 19234
rect 29486 19182 29538 19234
rect 30494 19182 30546 19234
rect 31502 19182 31554 19234
rect 32734 19182 32786 19234
rect 32958 19182 33010 19234
rect 33854 19182 33906 19234
rect 34302 19182 34354 19234
rect 34414 19182 34466 19234
rect 46622 19182 46674 19234
rect 46958 19182 47010 19234
rect 47630 19182 47682 19234
rect 50766 19182 50818 19234
rect 51326 19182 51378 19234
rect 51550 19182 51602 19234
rect 53230 19182 53282 19234
rect 53566 19182 53618 19234
rect 7422 19070 7474 19122
rect 9214 19070 9266 19122
rect 12126 19070 12178 19122
rect 13582 19070 13634 19122
rect 16046 19070 16098 19122
rect 19294 19070 19346 19122
rect 21534 19070 21586 19122
rect 27134 19070 27186 19122
rect 52894 19070 52946 19122
rect 1710 18958 1762 19010
rect 8654 18958 8706 19010
rect 12910 18958 12962 19010
rect 20750 18958 20802 19010
rect 22766 18958 22818 19010
rect 23102 18958 23154 19010
rect 28030 18958 28082 19010
rect 32398 18958 32450 19010
rect 41806 18958 41858 19010
rect 46062 18958 46114 19010
rect 46286 18958 46338 19010
rect 47182 18958 47234 19010
rect 50542 18958 50594 19010
rect 50878 18958 50930 19010
rect 50990 18958 51042 19010
rect 53678 18958 53730 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 7870 18622 7922 18674
rect 8654 18622 8706 18674
rect 11006 18622 11058 18674
rect 18062 18622 18114 18674
rect 18174 18622 18226 18674
rect 24446 18622 24498 18674
rect 24558 18622 24610 18674
rect 29598 18622 29650 18674
rect 34526 18622 34578 18674
rect 39566 18622 39618 18674
rect 6750 18510 6802 18562
rect 13134 18510 13186 18562
rect 14478 18510 14530 18562
rect 15262 18510 15314 18562
rect 16942 18510 16994 18562
rect 17838 18510 17890 18562
rect 17950 18510 18002 18562
rect 19182 18510 19234 18562
rect 21198 18510 21250 18562
rect 25678 18510 25730 18562
rect 27694 18510 27746 18562
rect 28366 18510 28418 18562
rect 34414 18510 34466 18562
rect 35198 18510 35250 18562
rect 41246 18510 41298 18562
rect 42590 18510 42642 18562
rect 43374 18510 43426 18562
rect 45726 18510 45778 18562
rect 47070 18510 47122 18562
rect 51998 18510 52050 18562
rect 54238 18510 54290 18562
rect 55134 18510 55186 18562
rect 6974 18398 7026 18450
rect 7198 18398 7250 18450
rect 9102 18398 9154 18450
rect 11790 18398 11842 18450
rect 12350 18398 12402 18450
rect 12798 18398 12850 18450
rect 13694 18398 13746 18450
rect 14814 18398 14866 18450
rect 16046 18398 16098 18450
rect 17502 18398 17554 18450
rect 19070 18398 19122 18450
rect 20750 18398 20802 18450
rect 21758 18398 21810 18450
rect 23214 18398 23266 18450
rect 25454 18398 25506 18450
rect 26126 18398 26178 18450
rect 27582 18398 27634 18450
rect 28142 18398 28194 18450
rect 29038 18398 29090 18450
rect 30270 18398 30322 18450
rect 30382 18398 30434 18450
rect 30606 18398 30658 18450
rect 33182 18398 33234 18450
rect 33406 18398 33458 18450
rect 34750 18398 34802 18450
rect 35086 18398 35138 18450
rect 35758 18398 35810 18450
rect 37998 18398 38050 18450
rect 38334 18398 38386 18450
rect 38670 18398 38722 18450
rect 39790 18398 39842 18450
rect 41022 18398 41074 18450
rect 42142 18398 42194 18450
rect 42926 18398 42978 18450
rect 43262 18398 43314 18450
rect 43598 18398 43650 18450
rect 43934 18398 43986 18450
rect 44158 18398 44210 18450
rect 44830 18398 44882 18450
rect 45614 18398 45666 18450
rect 46622 18398 46674 18450
rect 47182 18398 47234 18450
rect 47294 18398 47346 18450
rect 47742 18398 47794 18450
rect 48974 18398 49026 18450
rect 49870 18398 49922 18450
rect 51102 18398 51154 18450
rect 52558 18398 52610 18450
rect 53790 18398 53842 18450
rect 55694 18398 55746 18450
rect 9662 18286 9714 18338
rect 10110 18286 10162 18338
rect 10558 18286 10610 18338
rect 11454 18286 11506 18338
rect 13806 18286 13858 18338
rect 18846 18286 18898 18338
rect 23662 18286 23714 18338
rect 26910 18286 26962 18338
rect 31054 18286 31106 18338
rect 31950 18286 32002 18338
rect 39230 18286 39282 18338
rect 45838 18286 45890 18338
rect 49198 18286 49250 18338
rect 50766 18286 50818 18338
rect 51550 18286 51602 18338
rect 7422 18174 7474 18226
rect 14702 18174 14754 18226
rect 24334 18174 24386 18226
rect 29822 18174 29874 18226
rect 32174 18174 32226 18226
rect 32510 18174 32562 18226
rect 33854 18174 33906 18226
rect 35198 18174 35250 18226
rect 41806 18174 41858 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 30494 17838 30546 17890
rect 34302 17838 34354 17890
rect 42814 17838 42866 17890
rect 45502 17838 45554 17890
rect 49198 17838 49250 17890
rect 49534 17838 49586 17890
rect 9998 17726 10050 17778
rect 11902 17726 11954 17778
rect 12910 17726 12962 17778
rect 27022 17726 27074 17778
rect 28142 17726 28194 17778
rect 30606 17726 30658 17778
rect 33742 17726 33794 17778
rect 36542 17726 36594 17778
rect 37550 17726 37602 17778
rect 46846 17726 46898 17778
rect 48974 17726 49026 17778
rect 52558 17726 52610 17778
rect 54350 17726 54402 17778
rect 57934 17726 57986 17778
rect 9550 17614 9602 17666
rect 10670 17614 10722 17666
rect 11342 17614 11394 17666
rect 12462 17614 12514 17666
rect 13918 17614 13970 17666
rect 14366 17614 14418 17666
rect 15822 17614 15874 17666
rect 16830 17614 16882 17666
rect 18286 17614 18338 17666
rect 18622 17614 18674 17666
rect 20414 17614 20466 17666
rect 21422 17614 21474 17666
rect 23774 17614 23826 17666
rect 24446 17614 24498 17666
rect 25118 17614 25170 17666
rect 29598 17614 29650 17666
rect 30718 17614 30770 17666
rect 33182 17614 33234 17666
rect 35086 17614 35138 17666
rect 37214 17614 37266 17666
rect 38782 17614 38834 17666
rect 39342 17614 39394 17666
rect 40910 17614 40962 17666
rect 41694 17614 41746 17666
rect 45502 17614 45554 17666
rect 46398 17614 46450 17666
rect 50430 17614 50482 17666
rect 50990 17614 51042 17666
rect 52670 17614 52722 17666
rect 54574 17614 54626 17666
rect 55582 17614 55634 17666
rect 17166 17502 17218 17554
rect 18174 17502 18226 17554
rect 21646 17502 21698 17554
rect 21982 17502 22034 17554
rect 22542 17502 22594 17554
rect 23438 17502 23490 17554
rect 24110 17502 24162 17554
rect 31950 17502 32002 17554
rect 34190 17502 34242 17554
rect 34750 17502 34802 17554
rect 34862 17502 34914 17554
rect 37774 17502 37826 17554
rect 37886 17502 37938 17554
rect 38222 17502 38274 17554
rect 38446 17502 38498 17554
rect 39006 17502 39058 17554
rect 41134 17502 41186 17554
rect 42590 17502 42642 17554
rect 42702 17502 42754 17554
rect 45166 17502 45218 17554
rect 51102 17502 51154 17554
rect 52894 17502 52946 17554
rect 53454 17502 53506 17554
rect 55134 17502 55186 17554
rect 1710 17390 1762 17442
rect 7982 17390 8034 17442
rect 8430 17390 8482 17442
rect 8878 17390 8930 17442
rect 9326 17390 9378 17442
rect 11118 17390 11170 17442
rect 13582 17390 13634 17442
rect 16270 17390 16322 17442
rect 20750 17390 20802 17442
rect 22990 17390 23042 17442
rect 24782 17390 24834 17442
rect 25230 17390 25282 17442
rect 25454 17390 25506 17442
rect 26126 17390 26178 17442
rect 26574 17390 26626 17442
rect 27582 17390 27634 17442
rect 28702 17390 28754 17442
rect 29374 17390 29426 17442
rect 31502 17390 31554 17442
rect 32510 17390 32562 17442
rect 32958 17390 33010 17442
rect 33630 17390 33682 17442
rect 33854 17390 33906 17442
rect 34302 17390 34354 17442
rect 35982 17390 36034 17442
rect 38894 17390 38946 17442
rect 39678 17390 39730 17442
rect 40126 17390 40178 17442
rect 42030 17390 42082 17442
rect 46734 17390 46786 17442
rect 46958 17390 47010 17442
rect 47294 17390 47346 17442
rect 47630 17390 47682 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 5406 17054 5458 17106
rect 7310 17054 7362 17106
rect 9886 17054 9938 17106
rect 17838 17054 17890 17106
rect 26910 17054 26962 17106
rect 27918 17054 27970 17106
rect 28142 17054 28194 17106
rect 32622 17054 32674 17106
rect 33070 17054 33122 17106
rect 33406 17054 33458 17106
rect 39678 17054 39730 17106
rect 39902 17054 39954 17106
rect 47070 17054 47122 17106
rect 53230 17054 53282 17106
rect 54350 17054 54402 17106
rect 54462 17054 54514 17106
rect 55246 17054 55298 17106
rect 6078 16942 6130 16994
rect 6526 16942 6578 16994
rect 7646 16942 7698 16994
rect 8990 16942 9042 16994
rect 10782 16942 10834 16994
rect 12014 16942 12066 16994
rect 23774 16942 23826 16994
rect 25902 16942 25954 16994
rect 34190 16942 34242 16994
rect 34414 16942 34466 16994
rect 34526 16942 34578 16994
rect 34974 16942 35026 16994
rect 35086 16942 35138 16994
rect 38222 16942 38274 16994
rect 41470 16942 41522 16994
rect 45054 16942 45106 16994
rect 46286 16942 46338 16994
rect 6974 16830 7026 16882
rect 8430 16830 8482 16882
rect 11566 16830 11618 16882
rect 13358 16830 13410 16882
rect 14030 16830 14082 16882
rect 15710 16830 15762 16882
rect 18174 16830 18226 16882
rect 18958 16830 19010 16882
rect 19854 16830 19906 16882
rect 20302 16830 20354 16882
rect 23214 16830 23266 16882
rect 24334 16830 24386 16882
rect 25566 16830 25618 16882
rect 26350 16830 26402 16882
rect 27470 16830 27522 16882
rect 27806 16830 27858 16882
rect 28366 16830 28418 16882
rect 29150 16830 29202 16882
rect 31390 16830 31442 16882
rect 33966 16830 34018 16882
rect 35310 16830 35362 16882
rect 37550 16830 37602 16882
rect 38334 16830 38386 16882
rect 39118 16830 39170 16882
rect 39566 16830 39618 16882
rect 41358 16830 41410 16882
rect 44606 16830 44658 16882
rect 45502 16830 45554 16882
rect 46734 16830 46786 16882
rect 53566 16830 53618 16882
rect 55022 16830 55074 16882
rect 5742 16718 5794 16770
rect 13806 16718 13858 16770
rect 16158 16718 16210 16770
rect 22430 16718 22482 16770
rect 23886 16718 23938 16770
rect 25678 16718 25730 16770
rect 29486 16718 29538 16770
rect 31838 16718 31890 16770
rect 36990 16718 37042 16770
rect 38782 16718 38834 16770
rect 41806 16718 41858 16770
rect 45278 16718 45330 16770
rect 46062 16718 46114 16770
rect 46398 16718 46450 16770
rect 53342 16718 53394 16770
rect 7758 16606 7810 16658
rect 10334 16606 10386 16658
rect 22766 16606 22818 16658
rect 24110 16606 24162 16658
rect 54238 16606 54290 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 7870 16270 7922 16322
rect 8206 16270 8258 16322
rect 9998 16270 10050 16322
rect 10222 16270 10274 16322
rect 20078 16270 20130 16322
rect 31390 16270 31442 16322
rect 37774 16270 37826 16322
rect 42366 16270 42418 16322
rect 45166 16270 45218 16322
rect 52110 16270 52162 16322
rect 5854 16158 5906 16210
rect 11566 16158 11618 16210
rect 12014 16158 12066 16210
rect 12574 16158 12626 16210
rect 12910 16158 12962 16210
rect 14142 16158 14194 16210
rect 21646 16158 21698 16210
rect 26574 16158 26626 16210
rect 27918 16158 27970 16210
rect 32958 16158 33010 16210
rect 34302 16158 34354 16210
rect 42142 16158 42194 16210
rect 47182 16158 47234 16210
rect 49534 16158 49586 16210
rect 51774 16158 51826 16210
rect 53006 16158 53058 16210
rect 53678 16158 53730 16210
rect 6414 16046 6466 16098
rect 7086 16046 7138 16098
rect 8542 16046 8594 16098
rect 9102 16046 9154 16098
rect 9886 16046 9938 16098
rect 13470 16046 13522 16098
rect 14590 16046 14642 16098
rect 15374 16046 15426 16098
rect 15822 16046 15874 16098
rect 18174 16046 18226 16098
rect 19182 16046 19234 16098
rect 19966 16046 20018 16098
rect 20526 16046 20578 16098
rect 21758 16046 21810 16098
rect 23214 16046 23266 16098
rect 24558 16046 24610 16098
rect 25006 16046 25058 16098
rect 26238 16046 26290 16098
rect 26910 16046 26962 16098
rect 27470 16046 27522 16098
rect 29822 16046 29874 16098
rect 30830 16046 30882 16098
rect 33406 16046 33458 16098
rect 33742 16046 33794 16098
rect 37774 16046 37826 16098
rect 39566 16046 39618 16098
rect 39902 16046 39954 16098
rect 41470 16046 41522 16098
rect 43934 16046 43986 16098
rect 45166 16046 45218 16098
rect 46174 16046 46226 16098
rect 46958 16046 47010 16098
rect 47518 16046 47570 16098
rect 47966 16046 48018 16098
rect 48190 16046 48242 16098
rect 51550 16046 51602 16098
rect 52894 16046 52946 16098
rect 6974 15934 7026 15986
rect 7646 15934 7698 15986
rect 14926 15934 14978 15986
rect 18398 15934 18450 15986
rect 22094 15934 22146 15986
rect 27582 15934 27634 15986
rect 30046 15934 30098 15986
rect 30942 15934 30994 15986
rect 37438 15934 37490 15986
rect 38558 15934 38610 15986
rect 44158 15934 44210 15986
rect 44830 15934 44882 15986
rect 47070 15934 47122 15986
rect 6078 15822 6130 15874
rect 6750 15822 6802 15874
rect 10670 15822 10722 15874
rect 18846 15822 18898 15874
rect 21310 15822 21362 15874
rect 21534 15822 21586 15874
rect 28590 15822 28642 15874
rect 36542 15822 36594 15874
rect 37102 15822 37154 15874
rect 39342 15822 39394 15874
rect 42702 15822 42754 15874
rect 48078 15822 48130 15874
rect 49646 15822 49698 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 10782 15486 10834 15538
rect 15822 15486 15874 15538
rect 23438 15486 23490 15538
rect 25342 15486 25394 15538
rect 26350 15486 26402 15538
rect 28814 15486 28866 15538
rect 33630 15486 33682 15538
rect 34638 15486 34690 15538
rect 35870 15486 35922 15538
rect 37102 15486 37154 15538
rect 37886 15486 37938 15538
rect 39790 15486 39842 15538
rect 51102 15486 51154 15538
rect 51214 15486 51266 15538
rect 52782 15486 52834 15538
rect 9550 15374 9602 15426
rect 10110 15374 10162 15426
rect 10446 15374 10498 15426
rect 11790 15374 11842 15426
rect 12686 15374 12738 15426
rect 16270 15374 16322 15426
rect 16830 15374 16882 15426
rect 19854 15374 19906 15426
rect 20414 15374 20466 15426
rect 21758 15374 21810 15426
rect 22542 15374 22594 15426
rect 25790 15374 25842 15426
rect 27358 15374 27410 15426
rect 28254 15374 28306 15426
rect 29150 15374 29202 15426
rect 30046 15374 30098 15426
rect 30158 15374 30210 15426
rect 31614 15374 31666 15426
rect 32062 15374 32114 15426
rect 33742 15374 33794 15426
rect 34302 15374 34354 15426
rect 34414 15374 34466 15426
rect 36430 15374 36482 15426
rect 38334 15374 38386 15426
rect 42030 15374 42082 15426
rect 43374 15374 43426 15426
rect 52670 15374 52722 15426
rect 5630 15262 5682 15314
rect 6526 15262 6578 15314
rect 8766 15262 8818 15314
rect 12462 15262 12514 15314
rect 12798 15262 12850 15314
rect 15262 15262 15314 15314
rect 16606 15262 16658 15314
rect 17614 15262 17666 15314
rect 17950 15262 18002 15314
rect 18510 15262 18562 15314
rect 19630 15262 19682 15314
rect 19966 15262 20018 15314
rect 20526 15262 20578 15314
rect 21422 15262 21474 15314
rect 22766 15262 22818 15314
rect 24334 15262 24386 15314
rect 25678 15262 25730 15314
rect 26798 15262 26850 15314
rect 27694 15262 27746 15314
rect 29374 15262 29426 15314
rect 30382 15262 30434 15314
rect 31166 15262 31218 15314
rect 31838 15262 31890 15314
rect 33182 15262 33234 15314
rect 33854 15262 33906 15314
rect 34974 15262 35026 15314
rect 36094 15262 36146 15314
rect 36990 15262 37042 15314
rect 38222 15262 38274 15314
rect 39230 15262 39282 15314
rect 42478 15262 42530 15314
rect 49086 15262 49138 15314
rect 49422 15262 49474 15314
rect 50542 15262 50594 15314
rect 50990 15262 51042 15314
rect 53566 15262 53618 15314
rect 6078 15150 6130 15202
rect 6638 15150 6690 15202
rect 14478 15150 14530 15202
rect 15038 15150 15090 15202
rect 18622 15150 18674 15202
rect 21758 15150 21810 15202
rect 24558 15150 24610 15202
rect 24670 15150 24722 15202
rect 32174 15150 32226 15202
rect 38670 15150 38722 15202
rect 40238 15150 40290 15202
rect 41246 15150 41298 15202
rect 42926 15150 42978 15202
rect 45950 15150 46002 15202
rect 48862 15150 48914 15202
rect 49758 15150 49810 15202
rect 49982 15150 50034 15202
rect 52894 15150 52946 15202
rect 53342 15150 53394 15202
rect 54238 15150 54290 15202
rect 8318 15038 8370 15090
rect 14702 15038 14754 15090
rect 18734 15038 18786 15090
rect 31278 15038 31330 15090
rect 50318 15038 50370 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 7646 14702 7698 14754
rect 25790 14702 25842 14754
rect 33294 14702 33346 14754
rect 37998 14702 38050 14754
rect 57934 14702 57986 14754
rect 7310 14590 7362 14642
rect 7534 14590 7586 14642
rect 8318 14590 8370 14642
rect 11342 14590 11394 14642
rect 11790 14590 11842 14642
rect 12798 14590 12850 14642
rect 14590 14590 14642 14642
rect 15374 14590 15426 14642
rect 16718 14590 16770 14642
rect 23774 14590 23826 14642
rect 26126 14590 26178 14642
rect 28590 14590 28642 14642
rect 33854 14590 33906 14642
rect 43598 14590 43650 14642
rect 45502 14590 45554 14642
rect 46398 14590 46450 14642
rect 49086 14590 49138 14642
rect 6190 14478 6242 14530
rect 6638 14478 6690 14530
rect 7758 14478 7810 14530
rect 8542 14478 8594 14530
rect 9214 14478 9266 14530
rect 9550 14478 9602 14530
rect 10222 14478 10274 14530
rect 11902 14478 11954 14530
rect 13022 14478 13074 14530
rect 13470 14478 13522 14530
rect 15934 14478 15986 14530
rect 18846 14478 18898 14530
rect 19406 14478 19458 14530
rect 19742 14478 19794 14530
rect 21198 14478 21250 14530
rect 21534 14478 21586 14530
rect 22318 14478 22370 14530
rect 22990 14478 23042 14530
rect 23998 14478 24050 14530
rect 24446 14478 24498 14530
rect 27470 14478 27522 14530
rect 29710 14478 29762 14530
rect 30158 14478 30210 14530
rect 31278 14478 31330 14530
rect 31950 14478 32002 14530
rect 32622 14478 32674 14530
rect 33630 14478 33682 14530
rect 33966 14478 34018 14530
rect 34190 14478 34242 14530
rect 36430 14478 36482 14530
rect 38670 14478 38722 14530
rect 40238 14478 40290 14530
rect 41022 14478 41074 14530
rect 41918 14478 41970 14530
rect 45390 14478 45442 14530
rect 46286 14478 46338 14530
rect 47182 14478 47234 14530
rect 47406 14478 47458 14530
rect 48750 14478 48802 14530
rect 50094 14478 50146 14530
rect 54238 14478 54290 14530
rect 55582 14478 55634 14530
rect 6414 14366 6466 14418
rect 9774 14366 9826 14418
rect 10446 14366 10498 14418
rect 10670 14366 10722 14418
rect 16270 14366 16322 14418
rect 19854 14366 19906 14418
rect 21422 14366 21474 14418
rect 21870 14366 21922 14418
rect 23662 14366 23714 14418
rect 24894 14366 24946 14418
rect 25454 14366 25506 14418
rect 26574 14366 26626 14418
rect 27134 14366 27186 14418
rect 27694 14366 27746 14418
rect 27918 14366 27970 14418
rect 34638 14366 34690 14418
rect 36094 14366 36146 14418
rect 36206 14366 36258 14418
rect 37102 14366 37154 14418
rect 37662 14366 37714 14418
rect 38894 14366 38946 14418
rect 40798 14366 40850 14418
rect 43150 14366 43202 14418
rect 45950 14366 46002 14418
rect 46734 14366 46786 14418
rect 47966 14366 48018 14418
rect 50878 14366 50930 14418
rect 54574 14366 54626 14418
rect 6974 14254 7026 14306
rect 9886 14254 9938 14306
rect 20190 14254 20242 14306
rect 22766 14254 22818 14306
rect 26014 14254 26066 14306
rect 28030 14254 28082 14306
rect 28254 14254 28306 14306
rect 29150 14254 29202 14306
rect 34974 14254 35026 14306
rect 35422 14254 35474 14306
rect 37886 14254 37938 14306
rect 42814 14254 42866 14306
rect 43486 14254 43538 14306
rect 46510 14254 46562 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 5966 13918 6018 13970
rect 11566 13918 11618 13970
rect 15486 13918 15538 13970
rect 24670 13918 24722 13970
rect 25678 13918 25730 13970
rect 30270 13918 30322 13970
rect 43486 13918 43538 13970
rect 10222 13806 10274 13858
rect 12014 13806 12066 13858
rect 14478 13806 14530 13858
rect 18174 13806 18226 13858
rect 25454 13806 25506 13858
rect 25902 13806 25954 13858
rect 30830 13806 30882 13858
rect 32510 13806 32562 13858
rect 41806 13806 41858 13858
rect 46062 13806 46114 13858
rect 51774 13806 51826 13858
rect 52222 13806 52274 13858
rect 7982 13694 8034 13746
rect 8430 13694 8482 13746
rect 9774 13694 9826 13746
rect 10670 13694 10722 13746
rect 11454 13694 11506 13746
rect 13246 13694 13298 13746
rect 14702 13694 14754 13746
rect 15598 13694 15650 13746
rect 16830 13694 16882 13746
rect 17838 13694 17890 13746
rect 18062 13694 18114 13746
rect 19518 13694 19570 13746
rect 20526 13694 20578 13746
rect 20974 13694 21026 13746
rect 23326 13694 23378 13746
rect 23550 13694 23602 13746
rect 27694 13694 27746 13746
rect 28366 13694 28418 13746
rect 28926 13694 28978 13746
rect 31054 13694 31106 13746
rect 32174 13694 32226 13746
rect 33742 13694 33794 13746
rect 34750 13694 34802 13746
rect 35534 13694 35586 13746
rect 36990 13694 37042 13746
rect 38446 13694 38498 13746
rect 39902 13694 39954 13746
rect 40014 13694 40066 13746
rect 43038 13694 43090 13746
rect 45390 13694 45442 13746
rect 51998 13694 52050 13746
rect 6526 13582 6578 13634
rect 7086 13582 7138 13634
rect 7534 13582 7586 13634
rect 8990 13582 9042 13634
rect 11118 13582 11170 13634
rect 16270 13582 16322 13634
rect 18734 13582 18786 13634
rect 21198 13582 21250 13634
rect 23774 13582 23826 13634
rect 25790 13582 25842 13634
rect 27582 13582 27634 13634
rect 31726 13582 31778 13634
rect 33182 13582 33234 13634
rect 37102 13582 37154 13634
rect 38894 13582 38946 13634
rect 41022 13582 41074 13634
rect 41694 13582 41746 13634
rect 45614 13582 45666 13634
rect 51886 13582 51938 13634
rect 7198 13470 7250 13522
rect 20414 13470 20466 13522
rect 23886 13470 23938 13522
rect 29262 13470 29314 13522
rect 37550 13470 37602 13522
rect 38670 13470 38722 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 14030 13134 14082 13186
rect 18286 13134 18338 13186
rect 32958 13134 33010 13186
rect 6750 13022 6802 13074
rect 12910 13022 12962 13074
rect 13806 13022 13858 13074
rect 15822 13022 15874 13074
rect 22654 13022 22706 13074
rect 25118 13022 25170 13074
rect 26238 13022 26290 13074
rect 31950 13022 32002 13074
rect 33742 13022 33794 13074
rect 35086 13022 35138 13074
rect 35870 13022 35922 13074
rect 37550 13022 37602 13074
rect 40910 13022 40962 13074
rect 41582 13022 41634 13074
rect 42366 13022 42418 13074
rect 43374 13022 43426 13074
rect 46958 13022 47010 13074
rect 52782 13022 52834 13074
rect 57934 13022 57986 13074
rect 6302 12910 6354 12962
rect 7086 12910 7138 12962
rect 8542 12910 8594 12962
rect 10222 12910 10274 12962
rect 12126 12910 12178 12962
rect 14366 12910 14418 12962
rect 15038 12910 15090 12962
rect 16942 12910 16994 12962
rect 17614 12910 17666 12962
rect 19070 12910 19122 12962
rect 19854 12910 19906 12962
rect 20638 12910 20690 12962
rect 21422 12910 21474 12962
rect 21870 12910 21922 12962
rect 22990 12910 23042 12962
rect 23998 12910 24050 12962
rect 25006 12910 25058 12962
rect 26126 12910 26178 12962
rect 26910 12910 26962 12962
rect 27358 12910 27410 12962
rect 28030 12910 28082 12962
rect 28366 12910 28418 12962
rect 28590 12910 28642 12962
rect 29262 12910 29314 12962
rect 30382 12910 30434 12962
rect 31390 12910 31442 12962
rect 32174 12910 32226 12962
rect 32510 12910 32562 12962
rect 33966 12910 34018 12962
rect 34302 12910 34354 12962
rect 37886 12910 37938 12962
rect 39006 12910 39058 12962
rect 39678 12910 39730 12962
rect 40686 12910 40738 12962
rect 43150 12910 43202 12962
rect 44270 12910 44322 12962
rect 46622 12910 46674 12962
rect 51326 12910 51378 12962
rect 51662 12910 51714 12962
rect 51774 12910 51826 12962
rect 53006 12910 53058 12962
rect 55918 12910 55970 12962
rect 7422 12798 7474 12850
rect 7870 12798 7922 12850
rect 9662 12798 9714 12850
rect 10110 12798 10162 12850
rect 19742 12798 19794 12850
rect 22318 12798 22370 12850
rect 22542 12798 22594 12850
rect 24222 12798 24274 12850
rect 24782 12798 24834 12850
rect 26238 12798 26290 12850
rect 33518 12798 33570 12850
rect 35534 12798 35586 12850
rect 37102 12798 37154 12850
rect 38446 12798 38498 12850
rect 41470 12798 41522 12850
rect 41918 12798 41970 12850
rect 43822 12798 43874 12850
rect 49758 12798 49810 12850
rect 50990 12798 51042 12850
rect 51102 12798 51154 12850
rect 52110 12798 52162 12850
rect 53678 12798 53730 12850
rect 8094 12686 8146 12738
rect 12350 12686 12402 12738
rect 20638 12686 20690 12738
rect 28142 12686 28194 12738
rect 28254 12686 28306 12738
rect 31390 12686 31442 12738
rect 35758 12686 35810 12738
rect 36318 12686 36370 12738
rect 38222 12686 38274 12738
rect 38558 12686 38610 12738
rect 41694 12686 41746 12738
rect 49422 12686 49474 12738
rect 51998 12686 52050 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 9102 12350 9154 12402
rect 9886 12350 9938 12402
rect 37774 12350 37826 12402
rect 38446 12350 38498 12402
rect 39342 12350 39394 12402
rect 39454 12350 39506 12402
rect 40126 12350 40178 12402
rect 42030 12350 42082 12402
rect 50430 12350 50482 12402
rect 51886 12350 51938 12402
rect 52334 12350 52386 12402
rect 55918 12350 55970 12402
rect 7310 12238 7362 12290
rect 11006 12238 11058 12290
rect 12462 12238 12514 12290
rect 13694 12238 13746 12290
rect 16270 12238 16322 12290
rect 26014 12238 26066 12290
rect 30382 12238 30434 12290
rect 33070 12238 33122 12290
rect 34078 12238 34130 12290
rect 35646 12238 35698 12290
rect 37326 12238 37378 12290
rect 40014 12238 40066 12290
rect 41246 12238 41298 12290
rect 43934 12238 43986 12290
rect 46174 12238 46226 12290
rect 48190 12238 48242 12290
rect 49086 12238 49138 12290
rect 49310 12238 49362 12290
rect 49982 12238 50034 12290
rect 51102 12238 51154 12290
rect 52670 12238 52722 12290
rect 53006 12238 53058 12290
rect 5854 12126 5906 12178
rect 6302 12126 6354 12178
rect 7534 12126 7586 12178
rect 7982 12126 8034 12178
rect 10334 12126 10386 12178
rect 10894 12126 10946 12178
rect 11566 12126 11618 12178
rect 12686 12126 12738 12178
rect 13246 12126 13298 12178
rect 13582 12126 13634 12178
rect 14590 12126 14642 12178
rect 14814 12126 14866 12178
rect 15934 12126 15986 12178
rect 16718 12126 16770 12178
rect 19070 12126 19122 12178
rect 19854 12126 19906 12178
rect 20750 12126 20802 12178
rect 21198 12126 21250 12178
rect 22766 12126 22818 12178
rect 24558 12126 24610 12178
rect 26238 12126 26290 12178
rect 27134 12126 27186 12178
rect 27358 12126 27410 12178
rect 29486 12126 29538 12178
rect 29822 12126 29874 12178
rect 30718 12126 30770 12178
rect 31614 12126 31666 12178
rect 33294 12126 33346 12178
rect 34526 12126 34578 12178
rect 35086 12126 35138 12178
rect 36430 12126 36482 12178
rect 37550 12126 37602 12178
rect 37886 12126 37938 12178
rect 38894 12126 38946 12178
rect 39566 12126 39618 12178
rect 42926 12126 42978 12178
rect 45054 12126 45106 12178
rect 45390 12126 45442 12178
rect 45726 12126 45778 12178
rect 46958 12126 47010 12178
rect 47518 12126 47570 12178
rect 48862 12126 48914 12178
rect 50206 12126 50258 12178
rect 50766 12126 50818 12178
rect 52110 12126 52162 12178
rect 52782 12126 52834 12178
rect 53454 12126 53506 12178
rect 54574 12126 54626 12178
rect 55246 12126 55298 12178
rect 55582 12126 55634 12178
rect 6862 12014 6914 12066
rect 11118 12014 11170 12066
rect 12574 12014 12626 12066
rect 14030 12014 14082 12066
rect 17726 12014 17778 12066
rect 18622 12014 18674 12066
rect 19742 12014 19794 12066
rect 23214 12014 23266 12066
rect 29710 12014 29762 12066
rect 31390 12014 31442 12066
rect 36878 12014 36930 12066
rect 47406 12014 47458 12066
rect 52222 12014 52274 12066
rect 54350 12014 54402 12066
rect 8318 11902 8370 11954
rect 14814 11902 14866 11954
rect 17390 11902 17442 11954
rect 17726 11902 17778 11954
rect 23326 11902 23378 11954
rect 24446 11902 24498 11954
rect 28366 11902 28418 11954
rect 31838 11902 31890 11954
rect 33406 11902 33458 11954
rect 40126 11902 40178 11954
rect 53230 11902 53282 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 7534 11454 7586 11506
rect 9774 11566 9826 11618
rect 8430 11454 8482 11506
rect 8654 11454 8706 11506
rect 8766 11454 8818 11506
rect 10670 11566 10722 11618
rect 20078 11566 20130 11618
rect 25118 11566 25170 11618
rect 30830 11566 30882 11618
rect 10110 11454 10162 11506
rect 10334 11454 10386 11506
rect 12574 11454 12626 11506
rect 14030 11454 14082 11506
rect 19070 11454 19122 11506
rect 21870 11454 21922 11506
rect 24446 11454 24498 11506
rect 27134 11454 27186 11506
rect 31390 11454 31442 11506
rect 38446 11454 38498 11506
rect 38894 11454 38946 11506
rect 39678 11566 39730 11618
rect 40238 11566 40290 11618
rect 40462 11566 40514 11618
rect 41246 11566 41298 11618
rect 42814 11566 42866 11618
rect 47182 11566 47234 11618
rect 48302 11566 48354 11618
rect 54350 11566 54402 11618
rect 39902 11454 39954 11506
rect 40238 11454 40290 11506
rect 41246 11454 41298 11506
rect 43598 11454 43650 11506
rect 46398 11454 46450 11506
rect 46734 11454 46786 11506
rect 53006 11454 53058 11506
rect 53902 11454 53954 11506
rect 11118 11342 11170 11394
rect 11566 11342 11618 11394
rect 12126 11342 12178 11394
rect 13694 11342 13746 11394
rect 14926 11342 14978 11394
rect 16270 11342 16322 11394
rect 16830 11342 16882 11394
rect 19182 11342 19234 11394
rect 19966 11342 20018 11394
rect 21310 11342 21362 11394
rect 23438 11342 23490 11394
rect 24334 11342 24386 11394
rect 26126 11342 26178 11394
rect 27246 11342 27298 11394
rect 27806 11342 27858 11394
rect 28254 11342 28306 11394
rect 29486 11342 29538 11394
rect 30830 11342 30882 11394
rect 31726 11342 31778 11394
rect 32398 11342 32450 11394
rect 34638 11342 34690 11394
rect 36318 11342 36370 11394
rect 37102 11342 37154 11394
rect 37550 11342 37602 11394
rect 37998 11342 38050 11394
rect 42030 11342 42082 11394
rect 42254 11342 42306 11394
rect 43374 11342 43426 11394
rect 46958 11342 47010 11394
rect 47630 11342 47682 11394
rect 47966 11342 48018 11394
rect 48190 11342 48242 11394
rect 49086 11342 49138 11394
rect 49310 11342 49362 11394
rect 49422 11342 49474 11394
rect 54238 11342 54290 11394
rect 10670 11230 10722 11282
rect 11678 11230 11730 11282
rect 17614 11230 17666 11282
rect 22990 11230 23042 11282
rect 27022 11230 27074 11282
rect 28366 11230 28418 11282
rect 29262 11230 29314 11282
rect 29374 11230 29426 11282
rect 30494 11230 30546 11282
rect 32062 11230 32114 11282
rect 32286 11230 32338 11282
rect 36430 11230 36482 11282
rect 38782 11230 38834 11282
rect 42590 11230 42642 11282
rect 44270 11230 44322 11282
rect 47854 11230 47906 11282
rect 52782 11230 52834 11282
rect 6638 11118 6690 11170
rect 6974 11118 7026 11170
rect 7982 11118 8034 11170
rect 9326 11118 9378 11170
rect 9662 11118 9714 11170
rect 18062 11118 18114 11170
rect 20750 11118 20802 11170
rect 29934 11118 29986 11170
rect 31838 11118 31890 11170
rect 36206 11118 36258 11170
rect 38334 11118 38386 11170
rect 38558 11118 38610 11170
rect 39342 11118 39394 11170
rect 40686 11118 40738 11170
rect 41918 11118 41970 11170
rect 49870 11118 49922 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 7086 10782 7138 10834
rect 8094 10782 8146 10834
rect 10110 10782 10162 10834
rect 13918 10782 13970 10834
rect 14478 10782 14530 10834
rect 17726 10782 17778 10834
rect 21646 10782 21698 10834
rect 24110 10782 24162 10834
rect 24222 10782 24274 10834
rect 27582 10782 27634 10834
rect 32398 10782 32450 10834
rect 35086 10782 35138 10834
rect 37214 10782 37266 10834
rect 41694 10782 41746 10834
rect 42814 10782 42866 10834
rect 43374 10782 43426 10834
rect 43598 10782 43650 10834
rect 45950 10782 46002 10834
rect 50094 10782 50146 10834
rect 50318 10782 50370 10834
rect 51998 10782 52050 10834
rect 53790 10782 53842 10834
rect 8542 10670 8594 10722
rect 10334 10670 10386 10722
rect 12910 10670 12962 10722
rect 20862 10670 20914 10722
rect 22990 10670 23042 10722
rect 25230 10670 25282 10722
rect 26014 10670 26066 10722
rect 28590 10670 28642 10722
rect 31614 10670 31666 10722
rect 34526 10670 34578 10722
rect 36206 10670 36258 10722
rect 38222 10670 38274 10722
rect 48190 10670 48242 10722
rect 53006 10670 53058 10722
rect 53566 10670 53618 10722
rect 5742 10558 5794 10610
rect 6526 10558 6578 10610
rect 7534 10558 7586 10610
rect 7758 10558 7810 10610
rect 12014 10558 12066 10610
rect 12350 10558 12402 10610
rect 15262 10558 15314 10610
rect 15598 10558 15650 10610
rect 15822 10558 15874 10610
rect 16718 10558 16770 10610
rect 17950 10558 18002 10610
rect 18174 10558 18226 10610
rect 18622 10558 18674 10610
rect 19182 10558 19234 10610
rect 19742 10558 19794 10610
rect 20974 10558 21026 10610
rect 22206 10558 22258 10610
rect 24334 10558 24386 10610
rect 24670 10558 24722 10610
rect 25454 10558 25506 10610
rect 26238 10558 26290 10610
rect 26686 10558 26738 10610
rect 28814 10558 28866 10610
rect 29822 10558 29874 10610
rect 30270 10558 30322 10610
rect 31390 10558 31442 10610
rect 32286 10558 32338 10610
rect 33406 10558 33458 10610
rect 34302 10558 34354 10610
rect 35646 10558 35698 10610
rect 37662 10558 37714 10610
rect 41246 10558 41298 10610
rect 43262 10558 43314 10610
rect 44830 10558 44882 10610
rect 45166 10558 45218 10610
rect 46734 10558 46786 10610
rect 47518 10558 47570 10610
rect 48078 10558 48130 10610
rect 49646 10558 49698 10610
rect 51102 10558 51154 10610
rect 51214 10558 51266 10610
rect 6190 10446 6242 10498
rect 15038 10446 15090 10498
rect 15486 10446 15538 10498
rect 16270 10446 16322 10498
rect 18062 10446 18114 10498
rect 28142 10446 28194 10498
rect 28702 10446 28754 10498
rect 30718 10446 30770 10498
rect 33854 10446 33906 10498
rect 42926 10446 42978 10498
rect 46398 10446 46450 10498
rect 50206 10446 50258 10498
rect 50766 10446 50818 10498
rect 52782 10446 52834 10498
rect 53118 10446 53170 10498
rect 53902 10446 53954 10498
rect 8654 10334 8706 10386
rect 19406 10334 19458 10386
rect 40910 10334 40962 10386
rect 41246 10334 41298 10386
rect 42590 10334 42642 10386
rect 45502 10334 45554 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 13694 9998 13746 10050
rect 16158 9998 16210 10050
rect 20414 9998 20466 10050
rect 22206 9998 22258 10050
rect 27358 9998 27410 10050
rect 28366 9998 28418 10050
rect 33406 9998 33458 10050
rect 46846 9998 46898 10050
rect 47070 9998 47122 10050
rect 50766 9998 50818 10050
rect 50990 9998 51042 10050
rect 5966 9886 6018 9938
rect 7870 9886 7922 9938
rect 9886 9886 9938 9938
rect 14702 9886 14754 9938
rect 20190 9886 20242 9938
rect 23102 9886 23154 9938
rect 24670 9886 24722 9938
rect 32958 9886 33010 9938
rect 34750 9886 34802 9938
rect 35758 9886 35810 9938
rect 37102 9886 37154 9938
rect 38558 9886 38610 9938
rect 41470 9886 41522 9938
rect 45838 9886 45890 9938
rect 48638 9886 48690 9938
rect 50542 9886 50594 9938
rect 51438 9886 51490 9938
rect 7758 9774 7810 9826
rect 9438 9774 9490 9826
rect 10558 9774 10610 9826
rect 12238 9774 12290 9826
rect 12910 9774 12962 9826
rect 13806 9774 13858 9826
rect 14366 9774 14418 9826
rect 16046 9774 16098 9826
rect 17390 9774 17442 9826
rect 18510 9774 18562 9826
rect 19630 9774 19682 9826
rect 20414 9774 20466 9826
rect 21758 9774 21810 9826
rect 22094 9774 22146 9826
rect 22654 9774 22706 9826
rect 23886 9774 23938 9826
rect 24222 9774 24274 9826
rect 25118 9774 25170 9826
rect 26238 9774 26290 9826
rect 26686 9774 26738 9826
rect 27022 9774 27074 9826
rect 27806 9774 27858 9826
rect 28030 9774 28082 9826
rect 28254 9774 28306 9826
rect 29598 9774 29650 9826
rect 29934 9774 29986 9826
rect 31390 9774 31442 9826
rect 32510 9774 32562 9826
rect 34302 9774 34354 9826
rect 37438 9774 37490 9826
rect 37998 9774 38050 9826
rect 39566 9774 39618 9826
rect 39902 9774 39954 9826
rect 40350 9774 40402 9826
rect 41806 9774 41858 9826
rect 42254 9774 42306 9826
rect 46622 9774 46674 9826
rect 47854 9774 47906 9826
rect 48414 9774 48466 9826
rect 11678 9662 11730 9714
rect 12686 9662 12738 9714
rect 17166 9662 17218 9714
rect 17726 9662 17778 9714
rect 18174 9662 18226 9714
rect 39342 9662 39394 9714
rect 40574 9662 40626 9714
rect 41022 9662 41074 9714
rect 41694 9662 41746 9714
rect 42814 9662 42866 9714
rect 48974 9662 49026 9714
rect 51662 9662 51714 9714
rect 51774 9662 51826 9714
rect 6414 9550 6466 9602
rect 6862 9550 6914 9602
rect 7310 9550 7362 9602
rect 12798 9550 12850 9602
rect 13694 9550 13746 9602
rect 35310 9550 35362 9602
rect 36206 9550 36258 9602
rect 39566 9550 39618 9602
rect 42926 9550 42978 9602
rect 43150 9550 43202 9602
rect 43486 9550 43538 9602
rect 47518 9550 47570 9602
rect 51998 9550 52050 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 6526 9214 6578 9266
rect 6862 9214 6914 9266
rect 9102 9214 9154 9266
rect 9550 9214 9602 9266
rect 10446 9214 10498 9266
rect 14926 9214 14978 9266
rect 17614 9214 17666 9266
rect 22654 9214 22706 9266
rect 22766 9214 22818 9266
rect 24110 9214 24162 9266
rect 27694 9214 27746 9266
rect 29598 9214 29650 9266
rect 34078 9214 34130 9266
rect 39118 9214 39170 9266
rect 39566 9214 39618 9266
rect 40238 9214 40290 9266
rect 44158 9214 44210 9266
rect 45614 9214 45666 9266
rect 1710 9102 1762 9154
rect 7870 9102 7922 9154
rect 8318 9102 8370 9154
rect 9886 9102 9938 9154
rect 10222 9102 10274 9154
rect 13694 9102 13746 9154
rect 14142 9102 14194 9154
rect 17838 9102 17890 9154
rect 20750 9102 20802 9154
rect 23326 9102 23378 9154
rect 25566 9102 25618 9154
rect 28030 9102 28082 9154
rect 31502 9102 31554 9154
rect 33182 9102 33234 9154
rect 35870 9102 35922 9154
rect 36990 9102 37042 9154
rect 38782 9102 38834 9154
rect 42030 9102 42082 9154
rect 44606 9102 44658 9154
rect 44830 9102 44882 9154
rect 48750 9102 48802 9154
rect 48862 9102 48914 9154
rect 54014 9102 54066 9154
rect 6190 8990 6242 9042
rect 7758 8990 7810 9042
rect 11230 8990 11282 9042
rect 11902 8990 11954 9042
rect 12574 8990 12626 9042
rect 13134 8990 13186 9042
rect 14590 8990 14642 9042
rect 14926 8990 14978 9042
rect 15934 8990 15986 9042
rect 16270 8990 16322 9042
rect 19518 8990 19570 9042
rect 21086 8990 21138 9042
rect 21870 8990 21922 9042
rect 23662 8990 23714 9042
rect 24110 8990 24162 9042
rect 25454 8990 25506 9042
rect 27134 8990 27186 9042
rect 28590 8990 28642 9042
rect 29822 8990 29874 9042
rect 31838 8990 31890 9042
rect 33070 8990 33122 9042
rect 34190 8990 34242 9042
rect 36318 8990 36370 9042
rect 36766 8990 36818 9042
rect 41246 8990 41298 9042
rect 49086 8990 49138 9042
rect 52670 8990 52722 9042
rect 53342 8990 53394 9042
rect 53678 8990 53730 9042
rect 7422 8878 7474 8930
rect 11006 8878 11058 8930
rect 11454 8878 11506 8930
rect 13358 8878 13410 8930
rect 16158 8878 16210 8930
rect 18174 8878 18226 8930
rect 20526 8878 20578 8930
rect 21422 8878 21474 8930
rect 25342 8878 25394 8930
rect 34638 8878 34690 8930
rect 38222 8878 38274 8930
rect 41134 8878 41186 8930
rect 42814 8878 42866 8930
rect 44718 8878 44770 8930
rect 52558 8878 52610 8930
rect 10558 8766 10610 8818
rect 16718 8766 16770 8818
rect 18062 8766 18114 8818
rect 19518 8766 19570 8818
rect 22542 8766 22594 8818
rect 43934 8766 43986 8818
rect 44270 8766 44322 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19294 8430 19346 8482
rect 19966 8430 20018 8482
rect 44942 8430 44994 8482
rect 6302 8318 6354 8370
rect 9550 8318 9602 8370
rect 11902 8318 11954 8370
rect 12798 8318 12850 8370
rect 14702 8318 14754 8370
rect 19070 8318 19122 8370
rect 20638 8318 20690 8370
rect 24894 8318 24946 8370
rect 28478 8318 28530 8370
rect 30942 8318 30994 8370
rect 37438 8318 37490 8370
rect 37998 8318 38050 8370
rect 41246 8318 41298 8370
rect 45278 8318 45330 8370
rect 57934 8318 57986 8370
rect 6750 8206 6802 8258
rect 7198 8206 7250 8258
rect 8430 8206 8482 8258
rect 8878 8206 8930 8258
rect 11230 8206 11282 8258
rect 12238 8206 12290 8258
rect 13022 8206 13074 8258
rect 13358 8206 13410 8258
rect 13694 8206 13746 8258
rect 14590 8206 14642 8258
rect 14926 8206 14978 8258
rect 16494 8206 16546 8258
rect 17726 8206 17778 8258
rect 18734 8206 18786 8258
rect 19518 8206 19570 8258
rect 21982 8206 22034 8258
rect 22542 8206 22594 8258
rect 23102 8206 23154 8258
rect 24222 8206 24274 8258
rect 25790 8206 25842 8258
rect 27694 8206 27746 8258
rect 28030 8206 28082 8258
rect 29374 8206 29426 8258
rect 29934 8206 29986 8258
rect 32398 8206 32450 8258
rect 33630 8206 33682 8258
rect 35646 8206 35698 8258
rect 37102 8206 37154 8258
rect 40350 8206 40402 8258
rect 40574 8206 40626 8258
rect 45054 8206 45106 8258
rect 47742 8206 47794 8258
rect 47854 8206 47906 8258
rect 47966 8206 48018 8258
rect 48638 8206 48690 8258
rect 48974 8206 49026 8258
rect 49310 8206 49362 8258
rect 55582 8206 55634 8258
rect 7646 8094 7698 8146
rect 13582 8094 13634 8146
rect 14478 8094 14530 8146
rect 16382 8094 16434 8146
rect 20190 8094 20242 8146
rect 21646 8094 21698 8146
rect 24558 8094 24610 8146
rect 26350 8094 26402 8146
rect 28142 8094 28194 8146
rect 30606 8094 30658 8146
rect 30830 8094 30882 8146
rect 31950 8094 32002 8146
rect 34078 8094 34130 8146
rect 36318 8094 36370 8146
rect 37214 8094 37266 8146
rect 37550 8094 37602 8146
rect 38446 8094 38498 8146
rect 45390 8094 45442 8146
rect 45726 8094 45778 8146
rect 45950 8094 46002 8146
rect 46286 8094 46338 8146
rect 8206 7982 8258 8034
rect 9886 7982 9938 8034
rect 10334 7982 10386 8034
rect 10670 7982 10722 8034
rect 17614 7982 17666 8034
rect 26798 7982 26850 8034
rect 27246 7982 27298 8034
rect 30382 7982 30434 8034
rect 33406 7982 33458 8034
rect 34974 7982 35026 8034
rect 35870 7982 35922 8034
rect 46174 7982 46226 8034
rect 48414 7982 48466 8034
rect 48862 7982 48914 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 6862 7646 6914 7698
rect 7982 7646 8034 7698
rect 9102 7646 9154 7698
rect 15934 7646 15986 7698
rect 17614 7646 17666 7698
rect 17950 7646 18002 7698
rect 19070 7646 19122 7698
rect 20302 7646 20354 7698
rect 35086 7646 35138 7698
rect 36654 7646 36706 7698
rect 51550 7646 51602 7698
rect 12686 7534 12738 7586
rect 13806 7534 13858 7586
rect 15486 7534 15538 7586
rect 15710 7534 15762 7586
rect 16830 7534 16882 7586
rect 17838 7534 17890 7586
rect 20526 7534 20578 7586
rect 20638 7534 20690 7586
rect 23550 7534 23602 7586
rect 24670 7534 24722 7586
rect 25230 7534 25282 7586
rect 25342 7534 25394 7586
rect 26350 7534 26402 7586
rect 35534 7534 35586 7586
rect 38446 7534 38498 7586
rect 50654 7534 50706 7586
rect 9550 7422 9602 7474
rect 10110 7422 10162 7474
rect 11790 7422 11842 7474
rect 13358 7422 13410 7474
rect 13470 7422 13522 7474
rect 14142 7422 14194 7474
rect 15150 7422 15202 7474
rect 16046 7422 16098 7474
rect 17278 7422 17330 7474
rect 22094 7422 22146 7474
rect 22654 7422 22706 7474
rect 23214 7422 23266 7474
rect 24446 7422 24498 7474
rect 25902 7422 25954 7474
rect 27246 7422 27298 7474
rect 29150 7422 29202 7474
rect 30382 7422 30434 7474
rect 30830 7422 30882 7474
rect 31726 7422 31778 7474
rect 32286 7422 32338 7474
rect 33182 7422 33234 7474
rect 33742 7422 33794 7474
rect 34078 7422 34130 7474
rect 34302 7422 34354 7474
rect 34750 7422 34802 7474
rect 37326 7422 37378 7474
rect 37886 7422 37938 7474
rect 38670 7422 38722 7474
rect 39342 7422 39394 7474
rect 41134 7422 41186 7474
rect 43934 7422 43986 7474
rect 44606 7422 44658 7474
rect 45502 7422 45554 7474
rect 48862 7422 48914 7474
rect 48974 7422 49026 7474
rect 49310 7422 49362 7474
rect 50542 7422 50594 7474
rect 51438 7422 51490 7474
rect 7198 7310 7250 7362
rect 7758 7310 7810 7362
rect 8542 7310 8594 7362
rect 10782 7310 10834 7362
rect 11342 7310 11394 7362
rect 14702 7310 14754 7362
rect 18510 7310 18562 7362
rect 19742 7310 19794 7362
rect 21310 7310 21362 7362
rect 21758 7310 21810 7362
rect 23438 7310 23490 7362
rect 27806 7310 27858 7362
rect 29038 7310 29090 7362
rect 30718 7310 30770 7362
rect 34190 7310 34242 7362
rect 35646 7310 35698 7362
rect 36094 7310 36146 7362
rect 37998 7310 38050 7362
rect 39566 7310 39618 7362
rect 39678 7310 39730 7362
rect 40126 7310 40178 7362
rect 41582 7310 41634 7362
rect 46062 7310 46114 7362
rect 7198 7198 7250 7250
rect 7422 7198 7474 7250
rect 13694 7198 13746 7250
rect 18734 7198 18786 7250
rect 20638 7198 20690 7250
rect 25342 7198 25394 7250
rect 31950 7198 32002 7250
rect 35758 7198 35810 7250
rect 36318 7198 36370 7250
rect 38334 7198 38386 7250
rect 41918 7198 41970 7250
rect 49198 7198 49250 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 6862 6862 6914 6914
rect 7310 6862 7362 6914
rect 8206 6862 8258 6914
rect 14030 6862 14082 6914
rect 15598 6862 15650 6914
rect 35534 6862 35586 6914
rect 36542 6862 36594 6914
rect 45838 6862 45890 6914
rect 7310 6750 7362 6802
rect 7646 6750 7698 6802
rect 7982 6750 8034 6802
rect 15934 6750 15986 6802
rect 20190 6750 20242 6802
rect 22542 6750 22594 6802
rect 27806 6750 27858 6802
rect 29486 6750 29538 6802
rect 36206 6750 36258 6802
rect 37102 6750 37154 6802
rect 40798 6750 40850 6802
rect 45166 6750 45218 6802
rect 47742 6750 47794 6802
rect 50542 6750 50594 6802
rect 9326 6638 9378 6690
rect 10222 6638 10274 6690
rect 10782 6638 10834 6690
rect 11118 6638 11170 6690
rect 11790 6638 11842 6690
rect 12910 6638 12962 6690
rect 13582 6638 13634 6690
rect 14030 6638 14082 6690
rect 14926 6638 14978 6690
rect 16158 6638 16210 6690
rect 16606 6638 16658 6690
rect 17502 6638 17554 6690
rect 18398 6638 18450 6690
rect 18958 6638 19010 6690
rect 19294 6638 19346 6690
rect 19854 6638 19906 6690
rect 21422 6638 21474 6690
rect 22990 6638 23042 6690
rect 24670 6638 24722 6690
rect 26238 6638 26290 6690
rect 28254 6638 28306 6690
rect 29374 6638 29426 6690
rect 29934 6638 29986 6690
rect 30830 6638 30882 6690
rect 32286 6638 32338 6690
rect 34078 6638 34130 6690
rect 35198 6638 35250 6690
rect 37326 6638 37378 6690
rect 37998 6638 38050 6690
rect 40910 6638 40962 6690
rect 41358 6638 41410 6690
rect 42590 6638 42642 6690
rect 42814 6638 42866 6690
rect 43486 6638 43538 6690
rect 45278 6638 45330 6690
rect 49422 6638 49474 6690
rect 49870 6638 49922 6690
rect 50654 6638 50706 6690
rect 9886 6526 9938 6578
rect 16830 6526 16882 6578
rect 20078 6526 20130 6578
rect 21534 6526 21586 6578
rect 22094 6526 22146 6578
rect 22766 6526 22818 6578
rect 26126 6526 26178 6578
rect 28590 6526 28642 6578
rect 30606 6526 30658 6578
rect 34750 6526 34802 6578
rect 38446 6526 38498 6578
rect 41918 6526 41970 6578
rect 47966 6526 48018 6578
rect 51326 6526 51378 6578
rect 51662 6526 51714 6578
rect 8542 6414 8594 6466
rect 8990 6414 9042 6466
rect 15262 6414 15314 6466
rect 15822 6414 15874 6466
rect 16494 6414 16546 6466
rect 26686 6414 26738 6466
rect 27246 6414 27298 6466
rect 28478 6414 28530 6466
rect 34526 6414 34578 6466
rect 35646 6414 35698 6466
rect 39118 6414 39170 6466
rect 51998 6414 52050 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 7758 6078 7810 6130
rect 8094 6078 8146 6130
rect 8430 6078 8482 6130
rect 9774 6078 9826 6130
rect 11230 6078 11282 6130
rect 11678 6078 11730 6130
rect 12238 6078 12290 6130
rect 12798 6078 12850 6130
rect 16046 6078 16098 6130
rect 19406 6078 19458 6130
rect 26798 6078 26850 6130
rect 27806 6078 27858 6130
rect 35982 6078 36034 6130
rect 36542 6078 36594 6130
rect 37326 6078 37378 6130
rect 46734 6078 46786 6130
rect 47294 6078 47346 6130
rect 10670 5966 10722 6018
rect 14478 5966 14530 6018
rect 15262 5966 15314 6018
rect 18062 5966 18114 6018
rect 19182 5966 19234 6018
rect 24558 5966 24610 6018
rect 25230 5966 25282 6018
rect 27358 5966 27410 6018
rect 27582 5966 27634 6018
rect 30158 5966 30210 6018
rect 30606 5966 30658 6018
rect 32174 5966 32226 6018
rect 33630 5966 33682 6018
rect 35198 5966 35250 6018
rect 40238 5966 40290 6018
rect 46510 5966 46562 6018
rect 47182 5966 47234 6018
rect 10222 5854 10274 5906
rect 12574 5854 12626 5906
rect 13246 5854 13298 5906
rect 13694 5854 13746 5906
rect 13918 5854 13970 5906
rect 14254 5854 14306 5906
rect 14702 5854 14754 5906
rect 15038 5854 15090 5906
rect 17390 5854 17442 5906
rect 17838 5854 17890 5906
rect 19070 5854 19122 5906
rect 20190 5854 20242 5906
rect 21310 5854 21362 5906
rect 22206 5854 22258 5906
rect 23102 5854 23154 5906
rect 26238 5854 26290 5906
rect 28142 5854 28194 5906
rect 28814 5854 28866 5906
rect 29934 5854 29986 5906
rect 31166 5854 31218 5906
rect 31502 5854 31554 5906
rect 31950 5854 32002 5906
rect 32286 5854 32338 5906
rect 34078 5854 34130 5906
rect 34974 5854 35026 5906
rect 39790 5854 39842 5906
rect 40126 5854 40178 5906
rect 42030 5854 42082 5906
rect 42366 5854 42418 5906
rect 42590 5854 42642 5906
rect 47518 5854 47570 5906
rect 8990 5742 9042 5794
rect 14142 5742 14194 5794
rect 16382 5742 16434 5794
rect 16830 5742 16882 5794
rect 17614 5742 17666 5794
rect 18846 5742 18898 5794
rect 19742 5742 19794 5794
rect 27246 5742 27298 5794
rect 30046 5742 30098 5794
rect 30830 5742 30882 5794
rect 36878 5742 36930 5794
rect 46622 5742 46674 5794
rect 15374 5630 15426 5682
rect 15934 5630 15986 5682
rect 16382 5630 16434 5682
rect 23438 5630 23490 5682
rect 28254 5630 28306 5682
rect 39454 5630 39506 5682
rect 39790 5630 39842 5682
rect 58158 5630 58210 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 13470 5294 13522 5346
rect 16942 5294 16994 5346
rect 21422 5294 21474 5346
rect 27694 5294 27746 5346
rect 31614 5294 31666 5346
rect 9214 5182 9266 5234
rect 9662 5182 9714 5234
rect 10110 5182 10162 5234
rect 11566 5182 11618 5234
rect 13694 5182 13746 5234
rect 15150 5182 15202 5234
rect 16718 5182 16770 5234
rect 22542 5182 22594 5234
rect 24894 5182 24946 5234
rect 26574 5182 26626 5234
rect 27134 5182 27186 5234
rect 27358 5182 27410 5234
rect 28478 5182 28530 5234
rect 32062 5182 32114 5234
rect 33294 5182 33346 5234
rect 34302 5182 34354 5234
rect 35086 5182 35138 5234
rect 35422 5182 35474 5234
rect 38894 5182 38946 5234
rect 41134 5182 41186 5234
rect 45502 5182 45554 5234
rect 58158 5182 58210 5234
rect 10334 5070 10386 5122
rect 11118 5070 11170 5122
rect 12238 5070 12290 5122
rect 14030 5070 14082 5122
rect 14926 5070 14978 5122
rect 15374 5070 15426 5122
rect 15598 5070 15650 5122
rect 16270 5070 16322 5122
rect 16606 5070 16658 5122
rect 18286 5070 18338 5122
rect 19070 5070 19122 5122
rect 20302 5070 20354 5122
rect 20862 5070 20914 5122
rect 21310 5070 21362 5122
rect 22766 5070 22818 5122
rect 24446 5070 24498 5122
rect 26014 5070 26066 5122
rect 28142 5070 28194 5122
rect 29150 5070 29202 5122
rect 30830 5070 30882 5122
rect 32174 5070 32226 5122
rect 32398 5070 32450 5122
rect 33742 5070 33794 5122
rect 39342 5070 39394 5122
rect 39790 5070 39842 5122
rect 40126 5070 40178 5122
rect 40686 5070 40738 5122
rect 42814 5070 42866 5122
rect 43374 5070 43426 5122
rect 43486 5070 43538 5122
rect 43822 5070 43874 5122
rect 45166 5070 45218 5122
rect 46734 5070 46786 5122
rect 47406 5070 47458 5122
rect 48078 5070 48130 5122
rect 48638 5070 48690 5122
rect 10670 4958 10722 5010
rect 17502 4958 17554 5010
rect 18510 4958 18562 5010
rect 21422 4958 21474 5010
rect 26350 4958 26402 5010
rect 30046 4958 30098 5010
rect 41246 4958 41298 5010
rect 45390 4958 45442 5010
rect 46174 4958 46226 5010
rect 12574 4846 12626 4898
rect 13918 4846 13970 4898
rect 14142 4846 14194 4898
rect 14814 4846 14866 4898
rect 18062 4846 18114 4898
rect 18174 4846 18226 4898
rect 26462 4846 26514 4898
rect 26686 4846 26738 4898
rect 44158 4846 44210 4898
rect 48414 4846 48466 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 9774 4510 9826 4562
rect 10670 4510 10722 4562
rect 11230 4510 11282 4562
rect 13694 4510 13746 4562
rect 16046 4510 16098 4562
rect 17726 4510 17778 4562
rect 24782 4510 24834 4562
rect 27246 4510 27298 4562
rect 28366 4510 28418 4562
rect 29150 4510 29202 4562
rect 31614 4510 31666 4562
rect 33182 4510 33234 4562
rect 34190 4510 34242 4562
rect 34526 4510 34578 4562
rect 11902 4398 11954 4450
rect 12238 4398 12290 4450
rect 17614 4398 17666 4450
rect 17950 4398 18002 4450
rect 18846 4398 18898 4450
rect 25230 4398 25282 4450
rect 30942 4398 30994 4450
rect 40910 4398 40962 4450
rect 46286 4398 46338 4450
rect 58158 4398 58210 4450
rect 12910 4286 12962 4338
rect 13358 4286 13410 4338
rect 14254 4286 14306 4338
rect 14814 4286 14866 4338
rect 16270 4286 16322 4338
rect 18062 4286 18114 4338
rect 19294 4286 19346 4338
rect 19966 4286 20018 4338
rect 21534 4286 21586 4338
rect 21758 4286 21810 4338
rect 23438 4286 23490 4338
rect 25790 4286 25842 4338
rect 26462 4286 26514 4338
rect 27806 4286 27858 4338
rect 28590 4286 28642 4338
rect 29486 4286 29538 4338
rect 30606 4286 30658 4338
rect 31502 4286 31554 4338
rect 39678 4286 39730 4338
rect 40350 4286 40402 4338
rect 41134 4286 41186 4338
rect 47742 4286 47794 4338
rect 10334 4174 10386 4226
rect 11678 4174 11730 4226
rect 15262 4174 15314 4226
rect 16718 4174 16770 4226
rect 18958 4174 19010 4226
rect 20974 4174 21026 4226
rect 26798 4174 26850 4226
rect 29934 4174 29986 4226
rect 32174 4174 32226 4226
rect 33630 4174 33682 4226
rect 39902 4174 39954 4226
rect 46510 4174 46562 4226
rect 19182 4062 19234 4114
rect 22990 4062 23042 4114
rect 46622 4062 46674 4114
rect 47854 4062 47906 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 10334 3726 10386 3778
rect 12686 3726 12738 3778
rect 25790 3726 25842 3778
rect 26126 3726 26178 3778
rect 28590 3726 28642 3778
rect 29486 3726 29538 3778
rect 6974 3614 7026 3666
rect 10446 3614 10498 3666
rect 10894 3614 10946 3666
rect 11790 3614 11842 3666
rect 12238 3614 12290 3666
rect 12686 3614 12738 3666
rect 13358 3614 13410 3666
rect 13806 3614 13858 3666
rect 14142 3614 14194 3666
rect 16046 3614 16098 3666
rect 16494 3614 16546 3666
rect 17726 3614 17778 3666
rect 18510 3614 18562 3666
rect 18958 3614 19010 3666
rect 19406 3614 19458 3666
rect 20302 3614 20354 3666
rect 21310 3614 21362 3666
rect 21758 3614 21810 3666
rect 22094 3614 22146 3666
rect 23998 3614 24050 3666
rect 25118 3614 25170 3666
rect 27358 3614 27410 3666
rect 28590 3614 28642 3666
rect 29038 3614 29090 3666
rect 30158 3614 30210 3666
rect 30830 3614 30882 3666
rect 31278 3614 31330 3666
rect 33182 3614 33234 3666
rect 33630 3614 33682 3666
rect 34078 3614 34130 3666
rect 49086 3614 49138 3666
rect 52894 3614 52946 3666
rect 15598 3502 15650 3554
rect 17166 3502 17218 3554
rect 22430 3502 22482 3554
rect 23550 3502 23602 3554
rect 24558 3502 24610 3554
rect 26126 3502 26178 3554
rect 26686 3502 26738 3554
rect 27806 3502 27858 3554
rect 29710 3502 29762 3554
rect 31614 3502 31666 3554
rect 40910 3502 40962 3554
rect 44158 3502 44210 3554
rect 48414 3502 48466 3554
rect 52110 3502 52162 3554
rect 14590 3390 14642 3442
rect 15150 3390 15202 3442
rect 19854 3390 19906 3442
rect 23214 3390 23266 3442
rect 26462 3390 26514 3442
rect 29486 3390 29538 3442
rect 32398 3390 32450 3442
rect 4846 3278 4898 3330
rect 5630 3278 5682 3330
rect 7646 3278 7698 3330
rect 11342 3278 11394 3330
rect 32734 3278 32786 3330
rect 41470 3278 41522 3330
rect 44942 3278 44994 3330
rect 57710 3278 57762 3330
rect 58158 3278 58210 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 8064 59200 8176 60000
rect 10080 59200 10192 60000
rect 10752 59200 10864 60000
rect 13440 59200 13552 60000
rect 29568 59200 29680 60000
rect 47712 59200 47824 60000
rect 48384 59200 48496 60000
rect 49056 59200 49168 60000
rect 51072 59200 51184 60000
rect 52416 59200 52528 60000
rect 53088 59200 53200 60000
rect 53760 59200 53872 60000
rect 54432 59200 54544 60000
rect 55104 59200 55216 60000
rect 8092 55972 8148 59200
rect 10108 56308 10164 59200
rect 10332 56308 10388 56318
rect 10108 56306 10388 56308
rect 10108 56254 10334 56306
rect 10386 56254 10388 56306
rect 10108 56252 10388 56254
rect 10780 56308 10836 59200
rect 11004 56308 11060 56318
rect 10780 56306 11060 56308
rect 10780 56254 11006 56306
rect 11058 56254 11060 56306
rect 10780 56252 11060 56254
rect 13468 56308 13524 59200
rect 15372 57204 15428 57214
rect 13692 56308 13748 56318
rect 13468 56306 13748 56308
rect 13468 56254 13694 56306
rect 13746 56254 13748 56306
rect 13468 56252 13748 56254
rect 10332 56242 10388 56252
rect 11004 56242 11060 56252
rect 13692 56242 13748 56252
rect 8316 55972 8372 55982
rect 8092 55970 8372 55972
rect 8092 55918 8318 55970
rect 8370 55918 8372 55970
rect 8092 55916 8372 55918
rect 8316 55906 8372 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 1708 54626 1764 54638
rect 1708 54574 1710 54626
rect 1762 54574 1764 54626
rect 1708 53844 1764 54574
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 1708 53778 1764 53788
rect 14924 53508 14980 53518
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 14140 52276 14196 52286
rect 11900 51156 11956 51166
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 11228 49698 11284 49710
rect 11228 49646 11230 49698
rect 11282 49646 11284 49698
rect 11116 49586 11172 49598
rect 11116 49534 11118 49586
rect 11170 49534 11172 49586
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 8204 46564 8260 46574
rect 11116 46564 11172 49534
rect 11228 49588 11284 49646
rect 11228 48242 11284 49532
rect 11676 49700 11732 49710
rect 11676 49586 11732 49644
rect 11676 49534 11678 49586
rect 11730 49534 11732 49586
rect 11676 49522 11732 49534
rect 11676 48244 11732 48254
rect 11228 48190 11230 48242
rect 11282 48190 11284 48242
rect 11228 48178 11284 48190
rect 11340 48242 11732 48244
rect 11340 48190 11678 48242
rect 11730 48190 11732 48242
rect 11340 48188 11732 48190
rect 11228 46564 11284 46574
rect 11116 46508 11228 46564
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 8092 45220 8148 45230
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 1708 41300 1764 41310
rect 1708 41206 1764 41244
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 1708 37828 1764 37838
rect 1708 37734 1764 37772
rect 7868 37268 7924 37278
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 7868 35810 7924 37212
rect 7868 35758 7870 35810
rect 7922 35758 7924 35810
rect 7868 35746 7924 35758
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 8092 34692 8148 45164
rect 8092 34626 8148 34636
rect 4172 34132 4228 34142
rect 4172 34038 4228 34076
rect 4844 34132 4900 34142
rect 4844 34018 4900 34076
rect 4844 33966 4846 34018
rect 4898 33966 4900 34018
rect 1932 33908 1988 33918
rect 1932 33814 1988 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4844 33684 4900 33966
rect 4844 33618 4900 33628
rect 1932 33458 1988 33470
rect 1932 33406 1934 33458
rect 1986 33406 1988 33458
rect 1932 33012 1988 33406
rect 4284 33348 4340 33358
rect 4284 33254 4340 33292
rect 1932 32946 1988 32956
rect 1708 32674 1764 32686
rect 1708 32622 1710 32674
rect 1762 32622 1764 32674
rect 1708 32340 1764 32622
rect 1708 32274 1764 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 8204 31948 8260 46508
rect 11228 46470 11284 46508
rect 9884 46452 9940 46462
rect 9660 41970 9716 41982
rect 9660 41918 9662 41970
rect 9714 41918 9716 41970
rect 8876 41748 8932 41758
rect 8876 41298 8932 41692
rect 8876 41246 8878 41298
rect 8930 41246 8932 41298
rect 8876 41234 8932 41246
rect 9660 41188 9716 41918
rect 9884 41298 9940 46396
rect 10556 45332 10612 45342
rect 10108 44324 10164 44334
rect 9996 43540 10052 43550
rect 9996 41858 10052 43484
rect 10108 42866 10164 44268
rect 10332 44100 10388 44110
rect 10332 44006 10388 44044
rect 10444 43876 10500 43886
rect 10108 42814 10110 42866
rect 10162 42814 10164 42866
rect 10108 42802 10164 42814
rect 10220 43820 10444 43876
rect 10220 43538 10276 43820
rect 10444 43810 10500 43820
rect 10220 43486 10222 43538
rect 10274 43486 10276 43538
rect 9996 41806 9998 41858
rect 10050 41806 10052 41858
rect 9996 41794 10052 41806
rect 9884 41246 9886 41298
rect 9938 41246 9940 41298
rect 9884 41234 9940 41246
rect 10220 41300 10276 43486
rect 10444 43540 10500 43550
rect 10444 43446 10500 43484
rect 10220 41206 10276 41244
rect 10444 42754 10500 42766
rect 10444 42702 10446 42754
rect 10498 42702 10500 42754
rect 9436 41132 9660 41188
rect 8988 41074 9044 41086
rect 8988 41022 8990 41074
rect 9042 41022 9044 41074
rect 8764 40964 8820 40974
rect 8764 40870 8820 40908
rect 8988 40964 9044 41022
rect 9324 40964 9380 40974
rect 8988 40962 9380 40964
rect 8988 40910 9326 40962
rect 9378 40910 9380 40962
rect 8988 40908 9380 40910
rect 8540 39620 8596 39630
rect 8764 39620 8820 39630
rect 8540 39618 8764 39620
rect 8540 39566 8542 39618
rect 8594 39566 8764 39618
rect 8540 39564 8764 39566
rect 8540 39554 8596 39564
rect 8652 39058 8708 39564
rect 8764 39554 8820 39564
rect 8652 39006 8654 39058
rect 8706 39006 8708 39058
rect 8652 38994 8708 39006
rect 8764 38722 8820 38734
rect 8764 38670 8766 38722
rect 8818 38670 8820 38722
rect 8764 37828 8820 38670
rect 8988 38668 9044 40908
rect 9324 40898 9380 40908
rect 9436 40292 9492 41132
rect 9660 41122 9716 41132
rect 9772 40964 9828 40974
rect 9772 40404 9828 40908
rect 9100 40236 9604 40292
rect 9100 39730 9156 40236
rect 9100 39678 9102 39730
rect 9154 39678 9156 39730
rect 9100 39666 9156 39678
rect 9436 39620 9492 39630
rect 9436 39526 9492 39564
rect 8988 38612 9380 38668
rect 9100 37828 9156 37838
rect 8764 37826 9156 37828
rect 8764 37774 9102 37826
rect 9154 37774 9156 37826
rect 8764 37772 9156 37774
rect 8988 37604 9044 37614
rect 8988 37378 9044 37548
rect 8988 37326 8990 37378
rect 9042 37326 9044 37378
rect 8988 37314 9044 37326
rect 8316 37266 8372 37278
rect 8316 37214 8318 37266
rect 8370 37214 8372 37266
rect 8316 35812 8372 37214
rect 8316 35746 8372 35756
rect 8764 35698 8820 35710
rect 8764 35646 8766 35698
rect 8818 35646 8820 35698
rect 8764 34916 8820 35646
rect 8652 34914 8820 34916
rect 8652 34862 8766 34914
rect 8818 34862 8820 34914
rect 8652 34860 8820 34862
rect 8540 34244 8596 34254
rect 8652 34244 8708 34860
rect 8764 34850 8820 34860
rect 8988 34916 9044 34926
rect 8988 34822 9044 34860
rect 9100 34692 9156 37772
rect 9324 36372 9380 38612
rect 9548 37268 9604 40236
rect 9772 39732 9828 40348
rect 10220 40404 10276 40414
rect 10444 40404 10500 42702
rect 10556 40964 10612 45276
rect 10892 45218 10948 45230
rect 10892 45166 10894 45218
rect 10946 45166 10948 45218
rect 10892 44324 10948 45166
rect 11340 45108 11396 48188
rect 11676 48178 11732 48188
rect 11676 46676 11732 46686
rect 11228 45106 11396 45108
rect 11228 45054 11342 45106
rect 11394 45054 11396 45106
rect 11228 45052 11396 45054
rect 11452 46674 11732 46676
rect 11452 46622 11678 46674
rect 11730 46622 11732 46674
rect 11452 46620 11732 46622
rect 11452 45108 11508 46620
rect 11676 46610 11732 46620
rect 11900 46002 11956 51100
rect 12012 50708 12068 50718
rect 12012 49588 12068 50652
rect 12908 50708 12964 50718
rect 12908 50614 12964 50652
rect 13468 50708 13524 50718
rect 13468 50594 13524 50652
rect 13468 50542 13470 50594
rect 13522 50542 13524 50594
rect 13468 50530 13524 50542
rect 14140 50594 14196 52220
rect 14140 50542 14142 50594
rect 14194 50542 14196 50594
rect 14140 50530 14196 50542
rect 14364 51044 14420 51054
rect 13580 50370 13636 50382
rect 13580 50318 13582 50370
rect 13634 50318 13636 50370
rect 12460 49924 12516 49934
rect 12460 49922 13188 49924
rect 12460 49870 12462 49922
rect 12514 49870 13188 49922
rect 12460 49868 13188 49870
rect 12460 49858 12516 49868
rect 13132 49810 13188 49868
rect 13132 49758 13134 49810
rect 13186 49758 13188 49810
rect 13132 49746 13188 49758
rect 13580 49812 13636 50318
rect 13692 50372 13748 50382
rect 13692 50370 13972 50372
rect 13692 50318 13694 50370
rect 13746 50318 13972 50370
rect 13692 50316 13972 50318
rect 13692 50306 13748 50316
rect 13804 49812 13860 49822
rect 13580 49810 13860 49812
rect 13580 49758 13806 49810
rect 13858 49758 13860 49810
rect 13580 49756 13860 49758
rect 13804 49746 13860 49756
rect 12124 49700 12180 49710
rect 12124 49606 12180 49644
rect 12460 49700 12516 49710
rect 12012 49494 12068 49532
rect 12348 49588 12404 49598
rect 12460 49588 12516 49644
rect 13468 49700 13524 49710
rect 13468 49606 13524 49644
rect 12348 49586 12628 49588
rect 12348 49534 12350 49586
rect 12402 49534 12628 49586
rect 12348 49532 12628 49534
rect 12348 49522 12404 49532
rect 12348 47236 12404 47246
rect 12460 47236 12516 47246
rect 12348 47234 12460 47236
rect 12348 47182 12350 47234
rect 12402 47182 12460 47234
rect 12348 47180 12460 47182
rect 12348 47170 12404 47180
rect 11900 45950 11902 46002
rect 11954 45950 11956 46002
rect 11900 45938 11956 45950
rect 12348 46562 12404 46574
rect 12348 46510 12350 46562
rect 12402 46510 12404 46562
rect 12348 46116 12404 46510
rect 12460 46452 12516 47180
rect 12460 46386 12516 46396
rect 11564 45890 11620 45902
rect 11564 45838 11566 45890
rect 11618 45838 11620 45890
rect 11564 45332 11620 45838
rect 11564 45276 11956 45332
rect 11452 45052 11620 45108
rect 11116 44996 11172 45006
rect 11116 44902 11172 44940
rect 10780 44210 10836 44222
rect 10780 44158 10782 44210
rect 10834 44158 10836 44210
rect 10780 43540 10836 44158
rect 10780 43474 10836 43484
rect 10892 43538 10948 44268
rect 11228 43876 11284 45052
rect 11340 45042 11396 45052
rect 11228 43810 11284 43820
rect 11564 43764 11620 45052
rect 11900 45106 11956 45276
rect 11900 45054 11902 45106
rect 11954 45054 11956 45106
rect 11564 43708 11732 43764
rect 10892 43486 10894 43538
rect 10946 43486 10948 43538
rect 10892 43474 10948 43486
rect 11564 43538 11620 43550
rect 11564 43486 11566 43538
rect 11618 43486 11620 43538
rect 10892 43316 10948 43326
rect 10892 43222 10948 43260
rect 11004 43316 11060 43326
rect 11564 43316 11620 43486
rect 11004 43314 11564 43316
rect 11004 43262 11006 43314
rect 11058 43262 11564 43314
rect 11004 43260 11564 43262
rect 11004 43250 11060 43260
rect 11228 42866 11284 43260
rect 11564 43250 11620 43260
rect 11228 42814 11230 42866
rect 11282 42814 11284 42866
rect 11228 42802 11284 42814
rect 11676 42084 11732 43708
rect 11900 43426 11956 45054
rect 12236 44436 12292 44446
rect 12348 44436 12404 46060
rect 12460 46004 12516 46014
rect 12460 45910 12516 45948
rect 12236 44434 12404 44436
rect 12236 44382 12238 44434
rect 12290 44382 12404 44434
rect 12236 44380 12404 44382
rect 12236 44370 12292 44380
rect 11900 43374 11902 43426
rect 11954 43374 11956 43426
rect 11900 43362 11956 43374
rect 12012 44324 12068 44334
rect 11676 42028 11844 42084
rect 11564 41972 11620 41982
rect 11564 41970 11732 41972
rect 11564 41918 11566 41970
rect 11618 41918 11732 41970
rect 11564 41916 11732 41918
rect 11564 41906 11620 41916
rect 10780 41468 11396 41524
rect 10780 41186 10836 41468
rect 11004 41300 11060 41310
rect 11340 41300 11396 41468
rect 11060 41244 11172 41300
rect 11004 41234 11060 41244
rect 10780 41134 10782 41186
rect 10834 41134 10836 41186
rect 10780 41122 10836 41134
rect 10556 40908 10948 40964
rect 10668 40628 10724 40638
rect 10668 40514 10724 40572
rect 10668 40462 10670 40514
rect 10722 40462 10724 40514
rect 10668 40450 10724 40462
rect 10220 40402 10500 40404
rect 10220 40350 10222 40402
rect 10274 40350 10500 40402
rect 10220 40348 10500 40350
rect 10220 40338 10276 40348
rect 9884 39732 9940 39742
rect 9772 39730 9940 39732
rect 9772 39678 9886 39730
rect 9938 39678 9940 39730
rect 9772 39676 9940 39678
rect 9884 39666 9940 39676
rect 10332 38836 10388 40348
rect 10780 39396 10836 39406
rect 10332 38770 10388 38780
rect 10444 39394 10836 39396
rect 10444 39342 10782 39394
rect 10834 39342 10836 39394
rect 10444 39340 10836 39342
rect 10444 38834 10500 39340
rect 10780 39330 10836 39340
rect 10892 39172 10948 40908
rect 11116 40514 11172 41244
rect 11340 41298 11620 41300
rect 11340 41246 11342 41298
rect 11394 41246 11620 41298
rect 11340 41244 11620 41246
rect 11340 41234 11396 41244
rect 11116 40462 11118 40514
rect 11170 40462 11172 40514
rect 11116 40450 11172 40462
rect 11004 40404 11060 40414
rect 11004 40310 11060 40348
rect 11340 40404 11396 40414
rect 11340 39730 11396 40348
rect 11340 39678 11342 39730
rect 11394 39678 11396 39730
rect 11340 39666 11396 39678
rect 11564 39732 11620 41244
rect 10444 38782 10446 38834
rect 10498 38782 10500 38834
rect 9660 38050 9716 38062
rect 9660 37998 9662 38050
rect 9714 37998 9716 38050
rect 9660 37940 9716 37998
rect 9660 37874 9716 37884
rect 10444 37940 10500 38782
rect 10444 37874 10500 37884
rect 10780 39116 10948 39172
rect 11452 39396 11508 39406
rect 9660 37268 9716 37278
rect 9548 37266 9716 37268
rect 9548 37214 9662 37266
rect 9714 37214 9716 37266
rect 9548 37212 9716 37214
rect 9660 37156 9716 37212
rect 10556 37268 10612 37278
rect 10612 37212 10724 37268
rect 10556 37202 10612 37212
rect 9660 37090 9716 37100
rect 10108 36932 10164 36942
rect 9212 36260 9268 36270
rect 9212 36166 9268 36204
rect 9324 35138 9380 36316
rect 9996 36372 10052 36382
rect 9996 36278 10052 36316
rect 9548 35812 9604 35822
rect 9548 35718 9604 35756
rect 9324 35086 9326 35138
rect 9378 35086 9380 35138
rect 9324 35074 9380 35086
rect 9996 35698 10052 35710
rect 9996 35646 9998 35698
rect 10050 35646 10052 35698
rect 8596 34188 8708 34244
rect 8764 34636 9156 34692
rect 9996 34916 10052 35646
rect 8540 34018 8596 34188
rect 8540 33966 8542 34018
rect 8594 33966 8596 34018
rect 8540 33954 8596 33966
rect 1932 31892 1988 31902
rect 8204 31892 8372 31948
rect 1932 31798 1988 31836
rect 4284 31778 4340 31790
rect 4284 31726 4286 31778
rect 4338 31726 4340 31778
rect 4284 31556 4340 31726
rect 4732 31556 4788 31566
rect 4284 31554 4900 31556
rect 4284 31502 4734 31554
rect 4786 31502 4900 31554
rect 4284 31500 4900 31502
rect 4732 31490 4788 31500
rect 4284 30994 4340 31006
rect 4284 30942 4286 30994
rect 4338 30942 4340 30994
rect 1932 30884 1988 30894
rect 1932 30790 1988 30828
rect 4284 30436 4340 30942
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30370 4340 30380
rect 1708 30324 1764 30334
rect 1708 30230 1764 30268
rect 2156 29986 2212 29998
rect 2156 29934 2158 29986
rect 2210 29934 2212 29986
rect 2156 29652 2212 29934
rect 2156 29586 2212 29596
rect 4284 29540 4340 29550
rect 4284 29426 4340 29484
rect 4284 29374 4286 29426
rect 4338 29374 4340 29426
rect 4284 29362 4340 29374
rect 1932 29204 1988 29214
rect 4844 29204 4900 31500
rect 5628 30996 5684 31006
rect 6076 30996 6132 31006
rect 5628 30994 6020 30996
rect 5628 30942 5630 30994
rect 5682 30942 6020 30994
rect 5628 30940 6020 30942
rect 5628 30930 5684 30940
rect 4956 29204 5012 29214
rect 4844 29148 4956 29204
rect 1932 29110 1988 29148
rect 4956 29138 5012 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5964 28532 6020 30940
rect 6076 30902 6132 30940
rect 8316 29652 8372 31892
rect 8764 31668 8820 34636
rect 8988 34132 9044 34142
rect 9660 34132 9716 34142
rect 8988 34130 9940 34132
rect 8988 34078 8990 34130
rect 9042 34078 9662 34130
rect 9714 34078 9940 34130
rect 8988 34076 9940 34078
rect 8988 34066 9044 34076
rect 9660 34066 9716 34076
rect 8876 33348 8932 33358
rect 8876 32674 8932 33292
rect 8876 32622 8878 32674
rect 8930 32622 8932 32674
rect 8876 32564 8932 32622
rect 8876 32498 8932 32508
rect 9436 33122 9492 33134
rect 9436 33070 9438 33122
rect 9490 33070 9492 33122
rect 8988 32338 9044 32350
rect 8988 32286 8990 32338
rect 9042 32286 9044 32338
rect 8988 31780 9044 32286
rect 9436 31948 9492 33070
rect 9772 32562 9828 32574
rect 9772 32510 9774 32562
rect 9826 32510 9828 32562
rect 9772 31948 9828 32510
rect 8988 31714 9044 31724
rect 9100 31892 9828 31948
rect 8764 31602 8820 31612
rect 8540 31218 8596 31230
rect 8540 31166 8542 31218
rect 8594 31166 8596 31218
rect 8540 31108 8596 31166
rect 9100 31218 9156 31892
rect 9100 31166 9102 31218
rect 9154 31166 9156 31218
rect 9100 31154 9156 31166
rect 9884 31220 9940 34076
rect 9996 33348 10052 34860
rect 10108 34130 10164 36876
rect 10668 35924 10724 37212
rect 10780 36036 10836 39116
rect 11340 39060 11396 39070
rect 10892 38948 10948 38958
rect 10892 38854 10948 38892
rect 11340 38164 11396 39004
rect 11452 39058 11508 39340
rect 11452 39006 11454 39058
rect 11506 39006 11508 39058
rect 11452 38994 11508 39006
rect 11004 38108 11396 38164
rect 11004 38050 11060 38108
rect 11004 37998 11006 38050
rect 11058 37998 11060 38050
rect 11004 37986 11060 37998
rect 11116 37940 11172 37950
rect 10892 37268 10948 37278
rect 10892 37174 10948 37212
rect 11004 36482 11060 36494
rect 11004 36430 11006 36482
rect 11058 36430 11060 36482
rect 11004 36372 11060 36430
rect 11004 36306 11060 36316
rect 10780 35980 11060 36036
rect 10668 35868 10948 35924
rect 10780 35700 10836 35710
rect 10556 35698 10836 35700
rect 10556 35646 10782 35698
rect 10834 35646 10836 35698
rect 10556 35644 10836 35646
rect 10108 34078 10110 34130
rect 10162 34078 10164 34130
rect 10108 34066 10164 34078
rect 10444 34244 10500 34254
rect 10444 33570 10500 34188
rect 10444 33518 10446 33570
rect 10498 33518 10500 33570
rect 10444 33506 10500 33518
rect 9996 33254 10052 33292
rect 10556 33346 10612 35644
rect 10780 35634 10836 35644
rect 10892 35700 10948 35868
rect 10780 35028 10836 35038
rect 10780 34934 10836 34972
rect 10892 34914 10948 35644
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10892 34850 10948 34862
rect 10668 34244 10724 34254
rect 10668 34150 10724 34188
rect 10892 34132 10948 34142
rect 10556 33294 10558 33346
rect 10610 33294 10612 33346
rect 10556 33236 10612 33294
rect 10780 33348 10836 33358
rect 10892 33348 10948 34076
rect 10836 33292 10948 33348
rect 10780 33254 10836 33292
rect 10556 33170 10612 33180
rect 11004 33124 11060 35980
rect 11116 34130 11172 37884
rect 11228 37156 11284 37166
rect 11228 36594 11284 37100
rect 11228 36542 11230 36594
rect 11282 36542 11284 36594
rect 11228 36530 11284 36542
rect 11340 36036 11396 38108
rect 11452 38836 11508 38846
rect 11452 37938 11508 38780
rect 11452 37886 11454 37938
rect 11506 37886 11508 37938
rect 11452 36932 11508 37886
rect 11452 36866 11508 36876
rect 11452 36260 11508 36270
rect 11452 36166 11508 36204
rect 11228 35980 11396 36036
rect 11228 35588 11284 35980
rect 11340 35812 11396 35822
rect 11340 35718 11396 35756
rect 11228 35532 11396 35588
rect 11116 34078 11118 34130
rect 11170 34078 11172 34130
rect 11116 34066 11172 34078
rect 11228 33124 11284 33134
rect 11004 33122 11284 33124
rect 11004 33070 11230 33122
rect 11282 33070 11284 33122
rect 11004 33068 11284 33070
rect 10220 32564 10276 32574
rect 10220 32450 10276 32508
rect 10668 32564 10724 32574
rect 10668 32470 10724 32508
rect 10220 32398 10222 32450
rect 10274 32398 10276 32450
rect 10220 32386 10276 32398
rect 11116 32116 11172 33068
rect 11228 33058 11284 33068
rect 11228 32900 11284 32910
rect 11340 32900 11396 35532
rect 11284 32844 11396 32900
rect 11564 35028 11620 39676
rect 11676 39172 11732 41916
rect 11788 41524 11844 42028
rect 12012 42082 12068 44268
rect 12572 43988 12628 49532
rect 13804 49252 13860 49262
rect 13580 49138 13636 49150
rect 13580 49086 13582 49138
rect 13634 49086 13636 49138
rect 13580 49028 13636 49086
rect 13580 48962 13636 48972
rect 13356 48244 13412 48254
rect 13356 48150 13412 48188
rect 13804 48242 13860 49196
rect 13804 48190 13806 48242
rect 13858 48190 13860 48242
rect 13804 48178 13860 48190
rect 13916 48692 13972 50316
rect 14028 49588 14084 49598
rect 14028 49494 14084 49532
rect 13916 47570 13972 48636
rect 13916 47518 13918 47570
rect 13970 47518 13972 47570
rect 13916 47506 13972 47518
rect 14028 48802 14084 48814
rect 14028 48750 14030 48802
rect 14082 48750 14084 48802
rect 13580 47458 13636 47470
rect 13580 47406 13582 47458
rect 13634 47406 13636 47458
rect 13020 47234 13076 47246
rect 13020 47182 13022 47234
rect 13074 47182 13076 47234
rect 13020 46900 13076 47182
rect 13580 47012 13636 47406
rect 14028 47012 14084 48750
rect 13580 46946 13636 46956
rect 13916 46956 14084 47012
rect 14140 48244 14196 48254
rect 13020 46844 13524 46900
rect 13020 46676 13076 46686
rect 13468 46676 13524 46844
rect 13804 46676 13860 46686
rect 13020 46674 13412 46676
rect 13020 46622 13022 46674
rect 13074 46622 13412 46674
rect 13020 46620 13412 46622
rect 13468 46674 13860 46676
rect 13468 46622 13806 46674
rect 13858 46622 13860 46674
rect 13468 46620 13860 46622
rect 13020 46610 13076 46620
rect 12684 46452 12740 46462
rect 12684 46358 12740 46396
rect 13020 46452 13076 46462
rect 13020 46358 13076 46396
rect 13356 46116 13412 46620
rect 13692 46116 13748 46126
rect 13356 46060 13636 46116
rect 13468 45890 13524 45902
rect 13468 45838 13470 45890
rect 13522 45838 13524 45890
rect 12908 45668 12964 45678
rect 13468 45668 13524 45838
rect 12908 45666 13412 45668
rect 12908 45614 12910 45666
rect 12962 45614 13412 45666
rect 12908 45612 13412 45614
rect 12908 45602 12964 45612
rect 12796 45556 12852 45566
rect 12572 43922 12628 43932
rect 12684 45500 12796 45556
rect 12460 43650 12516 43662
rect 12460 43598 12462 43650
rect 12514 43598 12516 43650
rect 12012 42030 12014 42082
rect 12066 42030 12068 42082
rect 12012 42018 12068 42030
rect 12124 43538 12180 43550
rect 12124 43486 12126 43538
rect 12178 43486 12180 43538
rect 11788 41458 11844 41468
rect 11676 39106 11732 39116
rect 11788 41186 11844 41198
rect 11788 41134 11790 41186
rect 11842 41134 11844 41186
rect 11788 39618 11844 41134
rect 12012 40964 12068 41002
rect 12124 40964 12180 43486
rect 12460 43540 12516 43598
rect 12460 42532 12516 43484
rect 12460 42466 12516 42476
rect 12684 41748 12740 45500
rect 12796 45490 12852 45500
rect 13020 45106 13076 45118
rect 13020 45054 13022 45106
rect 13074 45054 13076 45106
rect 13020 44660 13076 45054
rect 13020 44594 13076 44604
rect 13356 43764 13412 45612
rect 13468 45602 13524 45612
rect 13580 43876 13636 46060
rect 13692 46022 13748 46060
rect 13692 44660 13748 44670
rect 13804 44660 13860 46620
rect 13748 44604 13860 44660
rect 13692 44594 13748 44604
rect 13916 44548 13972 46956
rect 14028 46788 14084 46798
rect 14140 46788 14196 48188
rect 14028 46786 14196 46788
rect 14028 46734 14030 46786
rect 14082 46734 14196 46786
rect 14028 46732 14196 46734
rect 14364 46786 14420 50988
rect 14588 50484 14644 50494
rect 14588 49476 14644 50428
rect 14812 50482 14868 50494
rect 14812 50430 14814 50482
rect 14866 50430 14868 50482
rect 14588 49410 14644 49420
rect 14700 49700 14756 49710
rect 14476 49364 14532 49374
rect 14476 49140 14532 49308
rect 14588 49140 14644 49150
rect 14476 49138 14644 49140
rect 14476 49086 14590 49138
rect 14642 49086 14644 49138
rect 14476 49084 14644 49086
rect 14364 46734 14366 46786
rect 14418 46734 14420 46786
rect 14028 46004 14084 46732
rect 14364 46722 14420 46734
rect 14028 45890 14084 45948
rect 14028 45838 14030 45890
rect 14082 45838 14084 45890
rect 14028 45826 14084 45838
rect 14140 46452 14196 46462
rect 14140 45890 14196 46396
rect 14588 46116 14644 49084
rect 14700 47236 14756 49644
rect 14812 49252 14868 50430
rect 14812 49186 14868 49196
rect 14700 47234 14868 47236
rect 14700 47182 14702 47234
rect 14754 47182 14868 47234
rect 14700 47180 14868 47182
rect 14700 47170 14756 47180
rect 14588 46050 14644 46060
rect 14700 46674 14756 46686
rect 14700 46622 14702 46674
rect 14754 46622 14756 46674
rect 14364 46004 14420 46014
rect 14140 45838 14142 45890
rect 14194 45838 14196 45890
rect 14140 45826 14196 45838
rect 14252 45892 14308 45902
rect 14252 45798 14308 45836
rect 14364 45890 14420 45948
rect 14364 45838 14366 45890
rect 14418 45838 14420 45890
rect 14364 45826 14420 45838
rect 14700 45780 14756 46622
rect 14588 45724 14756 45780
rect 14252 45668 14308 45678
rect 14140 44548 14196 44558
rect 13916 44492 14140 44548
rect 13580 43820 14084 43876
rect 13356 43708 13524 43764
rect 13020 43426 13076 43438
rect 13020 43374 13022 43426
rect 13074 43374 13076 43426
rect 13020 43316 13076 43374
rect 13020 42084 13076 43260
rect 13468 42756 13524 43708
rect 13580 43650 13636 43820
rect 13580 43598 13582 43650
rect 13634 43598 13636 43650
rect 13580 43586 13636 43598
rect 13692 43652 13748 43662
rect 13692 43650 13860 43652
rect 13692 43598 13694 43650
rect 13746 43598 13860 43650
rect 13692 43596 13860 43598
rect 13692 43586 13748 43596
rect 13692 43316 13748 43326
rect 13692 43222 13748 43260
rect 13468 42754 13748 42756
rect 13468 42702 13470 42754
rect 13522 42702 13748 42754
rect 13468 42700 13748 42702
rect 13468 42690 13524 42700
rect 13580 42532 13636 42542
rect 13244 42084 13300 42094
rect 13020 42028 13244 42084
rect 13244 41970 13300 42028
rect 13244 41918 13246 41970
rect 13298 41918 13300 41970
rect 13244 41906 13300 41918
rect 12684 41692 12852 41748
rect 12684 41524 12740 41534
rect 12348 41188 12404 41198
rect 12348 41094 12404 41132
rect 12684 41076 12740 41468
rect 12684 40982 12740 41020
rect 12068 40908 12180 40964
rect 12012 40898 12068 40908
rect 11788 39566 11790 39618
rect 11842 39566 11844 39618
rect 11788 38836 11844 39566
rect 12012 40740 12068 40750
rect 12012 39506 12068 40684
rect 12684 40292 12740 40302
rect 12684 39618 12740 40236
rect 12796 39730 12852 41692
rect 13468 41186 13524 41198
rect 13468 41134 13470 41186
rect 13522 41134 13524 41186
rect 13468 40740 13524 41134
rect 13580 41074 13636 42476
rect 13580 41022 13582 41074
rect 13634 41022 13636 41074
rect 13580 41010 13636 41022
rect 13468 40674 13524 40684
rect 13356 40628 13412 40638
rect 13244 40516 13300 40526
rect 13244 40422 13300 40460
rect 13356 40404 13412 40572
rect 13692 40404 13748 42700
rect 13804 41972 13860 43596
rect 13916 41972 13972 41982
rect 13804 41916 13916 41972
rect 13916 41878 13972 41916
rect 14028 41858 14084 43820
rect 14028 41806 14030 41858
rect 14082 41806 14084 41858
rect 14028 41748 14084 41806
rect 13356 40402 13524 40404
rect 13356 40350 13358 40402
rect 13410 40350 13524 40402
rect 13356 40348 13524 40350
rect 13356 40338 13412 40348
rect 13468 40292 13524 40348
rect 13468 40226 13524 40236
rect 13580 40402 13748 40404
rect 13580 40350 13694 40402
rect 13746 40350 13748 40402
rect 13580 40348 13748 40350
rect 12796 39678 12798 39730
rect 12850 39678 12852 39730
rect 12796 39666 12852 39678
rect 13580 39730 13636 40348
rect 13692 40338 13748 40348
rect 13916 41692 14084 41748
rect 13580 39678 13582 39730
rect 13634 39678 13636 39730
rect 12684 39566 12686 39618
rect 12738 39566 12740 39618
rect 12684 39554 12740 39566
rect 12908 39620 12964 39630
rect 12908 39526 12964 39564
rect 13580 39620 13636 39678
rect 13580 39554 13636 39564
rect 12012 39454 12014 39506
rect 12066 39454 12068 39506
rect 12012 39442 12068 39454
rect 12460 39396 12516 39406
rect 12460 39302 12516 39340
rect 13804 39396 13860 39406
rect 12124 38946 12180 38958
rect 12124 38894 12126 38946
rect 12178 38894 12180 38946
rect 11788 38770 11844 38780
rect 11900 38834 11956 38846
rect 11900 38782 11902 38834
rect 11954 38782 11956 38834
rect 11900 38724 11956 38782
rect 11900 38658 11956 38668
rect 12124 38668 12180 38894
rect 13468 38836 13524 38846
rect 13244 38724 13300 38762
rect 13468 38668 13524 38780
rect 12124 38612 12404 38668
rect 13244 38658 13300 38668
rect 12348 38050 12404 38612
rect 13356 38612 13524 38668
rect 12908 38164 12964 38174
rect 12908 38070 12964 38108
rect 12348 37998 12350 38050
rect 12402 37998 12404 38050
rect 12124 37938 12180 37950
rect 12124 37886 12126 37938
rect 12178 37886 12180 37938
rect 12124 37492 12180 37886
rect 12124 37426 12180 37436
rect 11676 35812 11732 35822
rect 11676 35718 11732 35756
rect 12348 35812 12404 37998
rect 12460 37380 12516 37390
rect 12460 37378 12628 37380
rect 12460 37326 12462 37378
rect 12514 37326 12628 37378
rect 12460 37324 12628 37326
rect 12460 37314 12516 37324
rect 12460 36594 12516 36606
rect 12460 36542 12462 36594
rect 12514 36542 12516 36594
rect 12460 36484 12516 36542
rect 12460 36418 12516 36428
rect 12348 35746 12404 35756
rect 12572 36372 12628 37324
rect 11900 35700 11956 35710
rect 11900 35606 11956 35644
rect 11228 32562 11284 32844
rect 11228 32510 11230 32562
rect 11282 32510 11284 32562
rect 11228 32498 11284 32510
rect 11116 32050 11172 32060
rect 11564 31948 11620 34972
rect 11788 35588 11844 35598
rect 11788 34914 11844 35532
rect 11788 34862 11790 34914
rect 11842 34862 11844 34914
rect 11788 34850 11844 34862
rect 12236 34804 12292 34814
rect 11676 34018 11732 34030
rect 11676 33966 11678 34018
rect 11730 33966 11732 34018
rect 11676 33684 11732 33966
rect 11676 33618 11732 33628
rect 12236 33458 12292 34748
rect 12572 34692 12628 36316
rect 12572 34626 12628 34636
rect 12796 37268 12852 37278
rect 12348 34132 12404 34142
rect 12348 34130 12740 34132
rect 12348 34078 12350 34130
rect 12402 34078 12740 34130
rect 12348 34076 12740 34078
rect 12348 34066 12404 34076
rect 12236 33406 12238 33458
rect 12290 33406 12292 33458
rect 12236 33394 12292 33406
rect 12684 33348 12740 34076
rect 12684 33254 12740 33292
rect 12124 33124 12180 33134
rect 10556 31892 10612 31902
rect 10556 31798 10612 31836
rect 11452 31892 11620 31948
rect 11788 32564 11844 32574
rect 11452 31890 11508 31892
rect 11452 31838 11454 31890
rect 11506 31838 11508 31890
rect 11452 31826 11508 31838
rect 9996 31780 10052 31790
rect 9996 31686 10052 31724
rect 10892 31780 10948 31790
rect 10892 31686 10948 31724
rect 11788 31778 11844 32508
rect 12124 32450 12180 33068
rect 12124 32398 12126 32450
rect 12178 32398 12180 32450
rect 12124 32386 12180 32398
rect 12460 32564 12516 32574
rect 12460 31948 12516 32508
rect 11788 31726 11790 31778
rect 11842 31726 11844 31778
rect 11788 31714 11844 31726
rect 12124 31892 12516 31948
rect 12796 32004 12852 37212
rect 12908 37044 12964 37054
rect 12908 36950 12964 36988
rect 13244 36372 13300 36382
rect 12908 36258 12964 36270
rect 12908 36206 12910 36258
rect 12962 36206 12964 36258
rect 12908 35252 12964 36206
rect 13244 35922 13300 36316
rect 13244 35870 13246 35922
rect 13298 35870 13300 35922
rect 13244 35858 13300 35870
rect 12908 35186 12964 35196
rect 12908 34914 12964 34926
rect 12908 34862 12910 34914
rect 12962 34862 12964 34914
rect 12908 34804 12964 34862
rect 12908 34738 12964 34748
rect 13356 33124 13412 38612
rect 13804 38052 13860 39340
rect 13804 37958 13860 37996
rect 13916 38164 13972 41692
rect 14028 39394 14084 39406
rect 14028 39342 14030 39394
rect 14082 39342 14084 39394
rect 14028 39060 14084 39342
rect 14028 38994 14084 39004
rect 13804 37268 13860 37278
rect 13916 37268 13972 38108
rect 14028 38052 14084 38062
rect 14028 37958 14084 37996
rect 13804 37266 13972 37268
rect 13804 37214 13806 37266
rect 13858 37214 13972 37266
rect 13804 37212 13972 37214
rect 13804 37202 13860 37212
rect 13692 37154 13748 37166
rect 14140 37156 14196 44492
rect 14252 42084 14308 45612
rect 14364 45332 14420 45342
rect 14364 45106 14420 45276
rect 14364 45054 14366 45106
rect 14418 45054 14420 45106
rect 14364 45042 14420 45054
rect 14476 44996 14532 45006
rect 14476 44902 14532 44940
rect 14588 44772 14644 45724
rect 14812 45668 14868 47180
rect 14924 46116 14980 53452
rect 15148 51378 15204 51390
rect 15148 51326 15150 51378
rect 15202 51326 15204 51378
rect 15148 50706 15204 51326
rect 15148 50654 15150 50706
rect 15202 50654 15204 50706
rect 15148 50642 15204 50654
rect 15036 50484 15092 50494
rect 15260 50484 15316 50522
rect 15036 50482 15204 50484
rect 15036 50430 15038 50482
rect 15090 50430 15204 50482
rect 15036 50428 15204 50430
rect 15036 50418 15092 50428
rect 15148 50372 15204 50428
rect 15260 50418 15316 50428
rect 15148 49812 15204 50316
rect 15260 49812 15316 49822
rect 15148 49756 15260 49812
rect 15260 49746 15316 49756
rect 15372 48468 15428 57148
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 25228 56308 25284 56318
rect 25228 56306 25844 56308
rect 25228 56254 25230 56306
rect 25282 56254 25844 56306
rect 25228 56252 25844 56254
rect 25228 56242 25284 56252
rect 25116 56082 25172 56094
rect 25116 56030 25118 56082
rect 25170 56030 25172 56082
rect 19180 55972 19236 55982
rect 19180 55970 19348 55972
rect 19180 55918 19182 55970
rect 19234 55918 19348 55970
rect 19180 55916 19348 55918
rect 19180 55906 19236 55916
rect 18060 55748 18116 55758
rect 17836 54740 17892 54750
rect 16828 53844 16884 53854
rect 16604 53842 16884 53844
rect 16604 53790 16830 53842
rect 16882 53790 16884 53842
rect 16604 53788 16884 53790
rect 16044 53620 16100 53630
rect 15596 52724 15652 52734
rect 15932 52724 15988 52734
rect 15596 52630 15652 52668
rect 15820 52722 15988 52724
rect 15820 52670 15934 52722
rect 15986 52670 15988 52722
rect 15820 52668 15988 52670
rect 15820 52274 15876 52668
rect 15932 52658 15988 52668
rect 15820 52222 15822 52274
rect 15874 52222 15876 52274
rect 15820 52210 15876 52222
rect 15484 51938 15540 51950
rect 15484 51886 15486 51938
rect 15538 51886 15540 51938
rect 15484 51604 15540 51886
rect 15484 51538 15540 51548
rect 15708 51938 15764 51950
rect 15708 51886 15710 51938
rect 15762 51886 15764 51938
rect 15484 51378 15540 51390
rect 15484 51326 15486 51378
rect 15538 51326 15540 51378
rect 15484 51268 15540 51326
rect 15484 51202 15540 51212
rect 15596 51266 15652 51278
rect 15596 51214 15598 51266
rect 15650 51214 15652 51266
rect 15484 50818 15540 50830
rect 15484 50766 15486 50818
rect 15538 50766 15540 50818
rect 15484 50428 15540 50766
rect 15596 50596 15652 51214
rect 15708 50932 15764 51886
rect 15932 51938 15988 51950
rect 15932 51886 15934 51938
rect 15986 51886 15988 51938
rect 15932 51380 15988 51886
rect 15708 50866 15764 50876
rect 15820 51378 15988 51380
rect 15820 51326 15934 51378
rect 15986 51326 15988 51378
rect 15820 51324 15988 51326
rect 16044 51380 16100 53564
rect 16492 53508 16548 53518
rect 16492 53414 16548 53452
rect 16604 53060 16660 53788
rect 16828 53778 16884 53788
rect 16940 53844 16996 53854
rect 16940 53730 16996 53788
rect 16940 53678 16942 53730
rect 16994 53678 16996 53730
rect 16940 53666 16996 53678
rect 17836 53844 17892 54684
rect 16716 53620 16772 53630
rect 16716 53526 16772 53564
rect 17836 53618 17892 53788
rect 17836 53566 17838 53618
rect 17890 53566 17892 53618
rect 17836 53554 17892 53566
rect 17164 53506 17220 53518
rect 17164 53454 17166 53506
rect 17218 53454 17220 53506
rect 17164 53284 17220 53454
rect 17500 53508 17556 53518
rect 17500 53414 17556 53452
rect 17164 53218 17220 53228
rect 17724 53172 17780 53182
rect 16380 53058 16660 53060
rect 16380 53006 16606 53058
rect 16658 53006 16660 53058
rect 16380 53004 16660 53006
rect 16380 52162 16436 53004
rect 16604 52994 16660 53004
rect 17500 53060 17556 53070
rect 16716 52948 16772 52958
rect 17276 52948 17332 52958
rect 16716 52946 17332 52948
rect 16716 52894 16718 52946
rect 16770 52894 17278 52946
rect 17330 52894 17332 52946
rect 16716 52892 17332 52894
rect 16716 52882 16772 52892
rect 17276 52882 17332 52892
rect 17500 52724 17556 53004
rect 17612 52948 17668 52958
rect 17612 52854 17668 52892
rect 17164 52668 17556 52724
rect 16940 52612 16996 52622
rect 16940 52164 16996 52556
rect 16380 52110 16382 52162
rect 16434 52110 16436 52162
rect 16380 52098 16436 52110
rect 16716 52162 16996 52164
rect 16716 52110 16942 52162
rect 16994 52110 16996 52162
rect 16716 52108 16996 52110
rect 16716 51940 16772 52108
rect 16940 52098 16996 52108
rect 16380 51884 16772 51940
rect 17164 52052 17220 52668
rect 16380 51492 16436 51884
rect 16716 51604 16772 51614
rect 16492 51492 16548 51502
rect 16380 51490 16548 51492
rect 16380 51438 16494 51490
rect 16546 51438 16548 51490
rect 16380 51436 16548 51438
rect 16268 51380 16324 51390
rect 16044 51324 16268 51380
rect 15596 50530 15652 50540
rect 15484 50372 15652 50428
rect 15260 48412 15428 48468
rect 15484 50260 15540 50270
rect 15036 46788 15092 46798
rect 15036 46694 15092 46732
rect 14924 46060 15092 46116
rect 14924 45892 14980 45902
rect 14924 45798 14980 45836
rect 14812 45602 14868 45612
rect 14924 45332 14980 45342
rect 15036 45332 15092 46060
rect 14980 45276 15092 45332
rect 14924 45266 14980 45276
rect 14476 44716 14644 44772
rect 15036 45106 15092 45118
rect 15036 45054 15038 45106
rect 15090 45054 15092 45106
rect 14364 44436 14420 44446
rect 14364 44342 14420 44380
rect 14252 42082 14420 42084
rect 14252 42030 14254 42082
rect 14306 42030 14420 42082
rect 14252 42028 14420 42030
rect 14252 42018 14308 42028
rect 14252 40402 14308 40414
rect 14252 40350 14254 40402
rect 14306 40350 14308 40402
rect 14252 40180 14308 40350
rect 14252 40114 14308 40124
rect 14364 39396 14420 42028
rect 14476 41748 14532 44716
rect 15036 44548 15092 45054
rect 15036 44482 15092 44492
rect 14588 44436 14644 44446
rect 14588 44322 14644 44380
rect 14588 44270 14590 44322
rect 14642 44270 14644 44322
rect 14588 44258 14644 44270
rect 14924 44324 14980 44334
rect 15148 44324 15204 44334
rect 14924 44322 15204 44324
rect 14924 44270 14926 44322
rect 14978 44270 15150 44322
rect 15202 44270 15204 44322
rect 14924 44268 15204 44270
rect 14924 44258 14980 44268
rect 15148 44258 15204 44268
rect 14700 44100 14756 44110
rect 14700 44098 14980 44100
rect 14700 44046 14702 44098
rect 14754 44046 14980 44098
rect 14700 44044 14980 44046
rect 14700 44034 14756 44044
rect 14588 43426 14644 43438
rect 14588 43374 14590 43426
rect 14642 43374 14644 43426
rect 14588 42084 14644 43374
rect 14588 42018 14644 42028
rect 14476 41682 14532 41692
rect 14812 41858 14868 41870
rect 14812 41806 14814 41858
rect 14866 41806 14868 41858
rect 14812 41412 14868 41806
rect 14812 41346 14868 41356
rect 14924 41860 14980 44044
rect 15036 42978 15092 42990
rect 15036 42926 15038 42978
rect 15090 42926 15092 42978
rect 15036 42084 15092 42926
rect 15260 42196 15316 48412
rect 15372 48242 15428 48254
rect 15372 48190 15374 48242
rect 15426 48190 15428 48242
rect 15372 48132 15428 48190
rect 15372 48066 15428 48076
rect 15484 48130 15540 50204
rect 15484 48078 15486 48130
rect 15538 48078 15540 48130
rect 15484 46788 15540 48078
rect 15596 47460 15652 50372
rect 15708 50372 15764 50382
rect 15708 50278 15764 50316
rect 15708 49698 15764 49710
rect 15708 49646 15710 49698
rect 15762 49646 15764 49698
rect 15708 48132 15764 49646
rect 15708 48066 15764 48076
rect 15596 47404 15764 47460
rect 15596 47236 15652 47246
rect 15596 47142 15652 47180
rect 15372 46732 15540 46788
rect 15372 45220 15428 46732
rect 15484 46564 15540 46574
rect 15484 46562 15652 46564
rect 15484 46510 15486 46562
rect 15538 46510 15652 46562
rect 15484 46508 15652 46510
rect 15484 46498 15540 46508
rect 15484 45890 15540 45902
rect 15484 45838 15486 45890
rect 15538 45838 15540 45890
rect 15484 45444 15540 45838
rect 15596 45892 15652 46508
rect 15596 45826 15652 45836
rect 15484 45378 15540 45388
rect 15596 45668 15652 45678
rect 15372 44436 15428 45164
rect 15372 44370 15428 44380
rect 15484 44098 15540 44110
rect 15484 44046 15486 44098
rect 15538 44046 15540 44098
rect 15484 43316 15540 44046
rect 15596 44100 15652 45612
rect 15708 44324 15764 47404
rect 15820 45892 15876 51324
rect 15932 51314 15988 51324
rect 16268 51286 16324 51324
rect 16380 51268 16436 51278
rect 16380 51174 16436 51212
rect 16380 50820 16436 50830
rect 16492 50820 16548 51436
rect 16380 50818 16548 50820
rect 16380 50766 16382 50818
rect 16434 50766 16548 50818
rect 16380 50764 16548 50766
rect 16716 51378 16772 51548
rect 16716 51326 16718 51378
rect 16770 51326 16772 51378
rect 16380 50754 16436 50764
rect 16380 50372 16436 50382
rect 16604 50372 16660 50382
rect 16380 50370 16660 50372
rect 16380 50318 16382 50370
rect 16434 50318 16606 50370
rect 16658 50318 16660 50370
rect 16380 50316 16660 50318
rect 16716 50372 16772 51326
rect 16940 50540 17108 50596
rect 16940 50482 16996 50540
rect 16940 50430 16942 50482
rect 16994 50430 16996 50482
rect 16940 50418 16996 50430
rect 17052 50484 17108 50540
rect 17164 50484 17220 51996
rect 17500 51268 17556 51278
rect 17500 51174 17556 51212
rect 17724 50820 17780 53116
rect 18060 52388 18116 55692
rect 19292 55188 19348 55916
rect 23772 55298 23828 55310
rect 23772 55246 23774 55298
rect 23826 55246 23828 55298
rect 19628 55188 19684 55198
rect 19292 55186 19684 55188
rect 19292 55134 19630 55186
rect 19682 55134 19684 55186
rect 19292 55132 19684 55134
rect 18732 55076 18788 55086
rect 18732 54740 18788 55020
rect 19180 55076 19236 55086
rect 19236 55020 19460 55076
rect 19180 54982 19236 55020
rect 18508 54684 18788 54740
rect 18508 53732 18564 54684
rect 19404 54626 19460 55020
rect 19404 54574 19406 54626
rect 19458 54574 19460 54626
rect 19404 54562 19460 54574
rect 18284 53676 18564 53732
rect 18620 54514 18676 54526
rect 18620 54462 18622 54514
rect 18674 54462 18676 54514
rect 18172 52612 18228 52622
rect 18284 52612 18340 53676
rect 18620 53284 18676 54462
rect 19068 54404 19124 54414
rect 19068 54310 19124 54348
rect 19292 53730 19348 53742
rect 19292 53678 19294 53730
rect 19346 53678 19348 53730
rect 18844 53284 18900 53294
rect 18620 53228 18844 53284
rect 18620 53060 18676 53070
rect 18620 52966 18676 53004
rect 18844 53058 18900 53228
rect 18844 53006 18846 53058
rect 18898 53006 18900 53058
rect 18228 52556 18340 52612
rect 18396 52946 18452 52958
rect 18396 52894 18398 52946
rect 18450 52894 18452 52946
rect 18396 52836 18452 52894
rect 18172 52546 18228 52556
rect 18060 52332 18228 52388
rect 17388 50818 17780 50820
rect 17388 50766 17726 50818
rect 17778 50766 17780 50818
rect 17388 50764 17780 50766
rect 17388 50708 17444 50764
rect 17724 50754 17780 50764
rect 18060 52164 18116 52174
rect 18060 50818 18116 52108
rect 18060 50766 18062 50818
rect 18114 50766 18116 50818
rect 18060 50754 18116 50766
rect 17388 50614 17444 50652
rect 17052 50428 17220 50484
rect 18172 50428 18228 52332
rect 18284 52276 18340 52286
rect 18396 52276 18452 52780
rect 18340 52220 18452 52276
rect 18508 52946 18564 52958
rect 18508 52894 18510 52946
rect 18562 52894 18564 52946
rect 18284 52210 18340 52220
rect 16716 50316 16884 50372
rect 16380 50260 16436 50316
rect 16604 50306 16660 50316
rect 15932 50204 16436 50260
rect 16828 50260 16884 50316
rect 16828 50204 16996 50260
rect 15932 46228 15988 50204
rect 16716 50148 16772 50158
rect 16268 49922 16324 49934
rect 16268 49870 16270 49922
rect 16322 49870 16324 49922
rect 16044 49812 16100 49822
rect 16044 49810 16212 49812
rect 16044 49758 16046 49810
rect 16098 49758 16212 49810
rect 16044 49756 16212 49758
rect 16044 49746 16100 49756
rect 16156 49026 16212 49756
rect 16156 48974 16158 49026
rect 16210 48974 16212 49026
rect 16156 48692 16212 48974
rect 16156 47460 16212 48636
rect 16268 48132 16324 49870
rect 16380 49922 16436 49934
rect 16380 49870 16382 49922
rect 16434 49870 16436 49922
rect 16380 49812 16436 49870
rect 16380 49746 16436 49756
rect 16716 49810 16772 50092
rect 16716 49758 16718 49810
rect 16770 49758 16772 49810
rect 16716 49746 16772 49758
rect 16828 49700 16884 49710
rect 16828 49606 16884 49644
rect 16940 49364 16996 50204
rect 17052 50148 17108 50158
rect 17164 50148 17220 50428
rect 17108 50092 17220 50148
rect 17948 50370 18004 50382
rect 17948 50318 17950 50370
rect 18002 50318 18004 50370
rect 17052 50082 17108 50092
rect 17836 49924 17892 49934
rect 17948 49924 18004 50318
rect 17892 49868 18004 49924
rect 18060 50372 18228 50428
rect 18284 51268 18340 51278
rect 17836 49830 17892 49868
rect 17500 49812 17556 49822
rect 17500 49718 17556 49756
rect 16940 49298 16996 49308
rect 17836 49364 17892 49374
rect 17836 49138 17892 49308
rect 17836 49086 17838 49138
rect 17890 49086 17892 49138
rect 17836 49074 17892 49086
rect 16604 49028 16660 49066
rect 17164 49028 17220 49038
rect 16604 48962 16660 48972
rect 17052 49026 17220 49028
rect 17052 48974 17166 49026
rect 17218 48974 17220 49026
rect 17052 48972 17220 48974
rect 16268 48038 16324 48076
rect 16604 48804 16660 48814
rect 16604 47682 16660 48748
rect 16604 47630 16606 47682
rect 16658 47630 16660 47682
rect 16604 47618 16660 47630
rect 16716 47570 16772 47582
rect 16716 47518 16718 47570
rect 16770 47518 16772 47570
rect 16268 47460 16324 47470
rect 16156 47458 16324 47460
rect 16156 47406 16270 47458
rect 16322 47406 16324 47458
rect 16156 47404 16324 47406
rect 16268 47394 16324 47404
rect 16716 47460 16772 47518
rect 16716 47394 16772 47404
rect 16044 47012 16100 47022
rect 16044 46898 16100 46956
rect 16044 46846 16046 46898
rect 16098 46846 16100 46898
rect 16044 46834 16100 46846
rect 16604 47012 16660 47022
rect 16268 46564 16324 46574
rect 16268 46470 16324 46508
rect 16492 46452 16548 46462
rect 15932 46172 16212 46228
rect 16044 46002 16100 46014
rect 16044 45950 16046 46002
rect 16098 45950 16100 46002
rect 15820 45836 15988 45892
rect 15820 44548 15876 44558
rect 15820 44454 15876 44492
rect 15932 44324 15988 45836
rect 16044 45780 16100 45950
rect 16044 45714 16100 45724
rect 15708 44268 15876 44324
rect 15708 44100 15764 44110
rect 15596 44098 15764 44100
rect 15596 44046 15710 44098
rect 15762 44046 15764 44098
rect 15596 44044 15764 44046
rect 15708 44034 15764 44044
rect 15708 43540 15764 43550
rect 15708 43446 15764 43484
rect 15820 43428 15876 44268
rect 15932 44230 15988 44268
rect 16156 43652 16212 46172
rect 16268 45892 16324 45902
rect 16268 45798 16324 45836
rect 16492 45556 16548 46396
rect 16604 45890 16660 46956
rect 16828 46900 16884 46910
rect 16828 46806 16884 46844
rect 16604 45838 16606 45890
rect 16658 45838 16660 45890
rect 16604 45826 16660 45838
rect 16716 46228 16772 46238
rect 16716 45778 16772 46172
rect 16828 46004 16884 46014
rect 16828 45892 16884 45948
rect 16940 45892 16996 45902
rect 16828 45836 16940 45892
rect 16940 45798 16996 45836
rect 16716 45726 16718 45778
rect 16770 45726 16772 45778
rect 16716 45714 16772 45726
rect 16492 45490 16548 45500
rect 16716 45220 16772 45230
rect 16772 45164 16996 45220
rect 16716 45126 16772 45164
rect 16268 45106 16324 45118
rect 16268 45054 16270 45106
rect 16322 45054 16324 45106
rect 16268 44996 16324 45054
rect 16268 44436 16324 44940
rect 16940 44884 16996 45164
rect 16268 44370 16324 44380
rect 16716 44436 16772 44446
rect 16380 44100 16436 44110
rect 16268 44098 16436 44100
rect 16268 44046 16382 44098
rect 16434 44046 16436 44098
rect 16268 44044 16436 44046
rect 16268 43764 16324 44044
rect 16380 44034 16436 44044
rect 16492 44100 16548 44110
rect 16492 44006 16548 44044
rect 16604 44098 16660 44110
rect 16604 44046 16606 44098
rect 16658 44046 16660 44098
rect 16268 43698 16324 43708
rect 16156 43586 16212 43596
rect 16380 43652 16436 43662
rect 16380 43558 16436 43596
rect 16604 43652 16660 44046
rect 16604 43586 16660 43596
rect 15820 43372 16212 43428
rect 15484 43092 15540 43260
rect 15484 43036 15876 43092
rect 15596 42868 15652 42878
rect 15260 42130 15316 42140
rect 15484 42866 15652 42868
rect 15484 42814 15598 42866
rect 15650 42814 15652 42866
rect 15484 42812 15652 42814
rect 15036 42018 15092 42028
rect 15260 41972 15316 41982
rect 15316 41916 15428 41972
rect 15260 41906 15316 41916
rect 15148 41860 15204 41870
rect 14924 41858 15204 41860
rect 14924 41806 15150 41858
rect 15202 41806 15204 41858
rect 14924 41804 15204 41806
rect 14924 41410 14980 41804
rect 15148 41794 15204 41804
rect 15260 41748 15316 41758
rect 15260 41654 15316 41692
rect 14924 41358 14926 41410
rect 14978 41358 14980 41410
rect 14924 41346 14980 41358
rect 15148 41636 15204 41646
rect 14588 41300 14644 41310
rect 14588 41186 14644 41244
rect 14588 41134 14590 41186
rect 14642 41134 14644 41186
rect 14588 41122 14644 41134
rect 14476 40962 14532 40974
rect 14476 40910 14478 40962
rect 14530 40910 14532 40962
rect 14476 40068 14532 40910
rect 15036 40962 15092 40974
rect 15036 40910 15038 40962
rect 15090 40910 15092 40962
rect 14812 40514 14868 40526
rect 14812 40462 14814 40514
rect 14866 40462 14868 40514
rect 14476 40002 14532 40012
rect 14700 40290 14756 40302
rect 14700 40238 14702 40290
rect 14754 40238 14756 40290
rect 14476 39732 14532 39742
rect 14532 39676 14644 39732
rect 14476 39638 14532 39676
rect 14364 39330 14420 39340
rect 14588 39058 14644 39676
rect 14588 39006 14590 39058
rect 14642 39006 14644 39058
rect 14588 38994 14644 39006
rect 14700 38388 14756 40238
rect 14812 40292 14868 40462
rect 15036 40404 15092 40910
rect 15148 40516 15204 41580
rect 15260 41300 15316 41310
rect 15260 41206 15316 41244
rect 15260 40628 15316 40638
rect 15372 40628 15428 41916
rect 15260 40626 15428 40628
rect 15260 40574 15262 40626
rect 15314 40574 15428 40626
rect 15260 40572 15428 40574
rect 15260 40562 15316 40572
rect 15148 40450 15204 40460
rect 15036 40292 15092 40348
rect 15036 40236 15204 40292
rect 14812 39060 14868 40236
rect 15148 39618 15204 40236
rect 15148 39566 15150 39618
rect 15202 39566 15204 39618
rect 15148 39554 15204 39566
rect 14812 38994 14868 39004
rect 15148 38948 15204 38958
rect 15148 38854 15204 38892
rect 14700 38322 14756 38332
rect 14476 38050 14532 38062
rect 14476 37998 14478 38050
rect 14530 37998 14532 38050
rect 13692 37102 13694 37154
rect 13746 37102 13748 37154
rect 13692 37044 13748 37102
rect 13916 37100 14196 37156
rect 14252 37380 14308 37390
rect 13916 37044 13972 37100
rect 13692 36988 13972 37044
rect 13804 36594 13860 36988
rect 13804 36542 13806 36594
rect 13858 36542 13860 36594
rect 13804 36530 13860 36542
rect 14140 36484 14196 36494
rect 14028 36370 14084 36382
rect 14028 36318 14030 36370
rect 14082 36318 14084 36370
rect 13692 35812 13748 35822
rect 13692 35698 13748 35756
rect 13692 35646 13694 35698
rect 13746 35646 13748 35698
rect 13692 35634 13748 35646
rect 14028 35588 14084 36318
rect 14140 35810 14196 36428
rect 14140 35758 14142 35810
rect 14194 35758 14196 35810
rect 14140 35746 14196 35758
rect 14028 35522 14084 35532
rect 14252 35364 14308 37324
rect 14028 35308 14308 35364
rect 14364 37042 14420 37054
rect 14364 36990 14366 37042
rect 14418 36990 14420 37042
rect 13356 33058 13412 33068
rect 13468 35252 13524 35262
rect 13468 32786 13524 35196
rect 14028 35026 14084 35308
rect 14028 34974 14030 35026
rect 14082 34974 14084 35026
rect 14028 34962 14084 34974
rect 13580 34692 13636 34702
rect 13636 34636 13748 34692
rect 13580 34598 13636 34636
rect 13580 34132 13636 34142
rect 13580 34038 13636 34076
rect 13692 33796 13748 34636
rect 13692 33730 13748 33740
rect 13468 32734 13470 32786
rect 13522 32734 13524 32786
rect 13468 32452 13524 32734
rect 14252 33236 14308 33246
rect 13468 32386 13524 32396
rect 13580 32676 13636 32686
rect 13580 31948 13636 32620
rect 14252 32674 14308 33180
rect 14252 32622 14254 32674
rect 14306 32622 14308 32674
rect 14028 32564 14084 32574
rect 14028 32470 14084 32508
rect 12796 31938 12852 31948
rect 13356 31892 13636 31948
rect 14140 32452 14196 32462
rect 12124 31666 12180 31892
rect 12124 31614 12126 31666
rect 12178 31614 12180 31666
rect 12124 31602 12180 31614
rect 9884 31154 9940 31164
rect 12348 31220 12404 31230
rect 12348 31126 12404 31164
rect 13356 31218 13412 31892
rect 14140 31778 14196 32396
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 14140 31714 14196 31726
rect 13356 31166 13358 31218
rect 13410 31166 13412 31218
rect 13356 31154 13412 31166
rect 14252 31220 14308 32622
rect 14364 31556 14420 36990
rect 14476 34690 14532 37998
rect 14924 36484 14980 36494
rect 14924 36482 15092 36484
rect 14924 36430 14926 36482
rect 14978 36430 15092 36482
rect 14924 36428 15092 36430
rect 14924 36418 14980 36428
rect 14588 35924 14644 35962
rect 14588 35858 14644 35868
rect 14588 35698 14644 35710
rect 14588 35646 14590 35698
rect 14642 35646 14644 35698
rect 14588 35588 14644 35646
rect 14588 35522 14644 35532
rect 14700 35252 14756 35262
rect 14756 35196 14868 35252
rect 14700 35186 14756 35196
rect 14476 34638 14478 34690
rect 14530 34638 14532 34690
rect 14476 33460 14532 34638
rect 14812 34914 14868 35196
rect 14812 34862 14814 34914
rect 14866 34862 14868 34914
rect 14700 34242 14756 34254
rect 14700 34190 14702 34242
rect 14754 34190 14756 34242
rect 14476 33394 14532 33404
rect 14588 34130 14644 34142
rect 14588 34078 14590 34130
rect 14642 34078 14644 34130
rect 14588 33908 14644 34078
rect 14588 32564 14644 33852
rect 14700 33236 14756 34190
rect 14812 33458 14868 34862
rect 14924 34916 14980 34926
rect 14924 34354 14980 34860
rect 15036 34804 15092 36428
rect 15036 34738 15092 34748
rect 15260 35698 15316 35710
rect 15260 35646 15262 35698
rect 15314 35646 15316 35698
rect 14924 34302 14926 34354
rect 14978 34302 14980 34354
rect 14924 34290 14980 34302
rect 15260 34356 15316 35646
rect 15372 35026 15428 40572
rect 15484 40626 15540 42812
rect 15596 42802 15652 42812
rect 15708 42754 15764 42766
rect 15708 42702 15710 42754
rect 15762 42702 15764 42754
rect 15596 42644 15652 42654
rect 15596 42194 15652 42588
rect 15596 42142 15598 42194
rect 15650 42142 15652 42194
rect 15596 42130 15652 42142
rect 15708 41972 15764 42702
rect 15820 42082 15876 43036
rect 16156 42420 16212 43372
rect 16380 43316 16436 43326
rect 16156 42364 16324 42420
rect 15820 42030 15822 42082
rect 15874 42030 15876 42082
rect 15820 42018 15876 42030
rect 16156 42196 16212 42206
rect 15708 41906 15764 41916
rect 16044 41972 16100 41982
rect 16044 41878 16100 41916
rect 16156 41858 16212 42140
rect 16156 41806 16158 41858
rect 16210 41806 16212 41858
rect 16156 41794 16212 41806
rect 16156 41524 16212 41534
rect 16044 41468 16156 41524
rect 15484 40574 15486 40626
rect 15538 40574 15540 40626
rect 15484 40404 15540 40574
rect 15708 40740 15764 40750
rect 15708 40626 15764 40684
rect 15708 40574 15710 40626
rect 15762 40574 15764 40626
rect 15708 40562 15764 40574
rect 15484 40338 15540 40348
rect 15596 40292 15652 40302
rect 15596 40198 15652 40236
rect 16044 39284 16100 41468
rect 16156 41458 16212 41468
rect 16268 41300 16324 42364
rect 16156 41298 16324 41300
rect 16156 41246 16270 41298
rect 16322 41246 16324 41298
rect 16156 41244 16324 41246
rect 16156 39396 16212 41244
rect 16268 41234 16324 41244
rect 16268 40516 16324 40526
rect 16268 40422 16324 40460
rect 16380 40292 16436 43260
rect 16604 42868 16660 42878
rect 16716 42868 16772 44380
rect 16940 44322 16996 44828
rect 17052 44548 17108 48972
rect 17164 48962 17220 48972
rect 17052 44482 17108 44492
rect 17164 48132 17220 48142
rect 16940 44270 16942 44322
rect 16994 44270 16996 44322
rect 16940 44258 16996 44270
rect 17052 44324 17108 44334
rect 17052 44210 17108 44268
rect 17052 44158 17054 44210
rect 17106 44158 17108 44210
rect 17052 44146 17108 44158
rect 17164 43708 17220 48076
rect 18060 48020 18116 50372
rect 18284 49140 18340 51212
rect 18396 51266 18452 51278
rect 18396 51214 18398 51266
rect 18450 51214 18452 51266
rect 18396 51156 18452 51214
rect 18396 51090 18452 51100
rect 18396 50820 18452 50830
rect 18508 50820 18564 52894
rect 18844 51380 18900 53006
rect 19292 53172 19348 53678
rect 19628 53732 19684 55132
rect 19964 55188 20020 55198
rect 19852 55076 19908 55114
rect 19964 55094 20020 55132
rect 20188 55186 20244 55198
rect 20188 55134 20190 55186
rect 20242 55134 20244 55186
rect 19852 55010 19908 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54516 20244 55134
rect 20860 55074 20916 55086
rect 21308 55076 21364 55086
rect 20860 55022 20862 55074
rect 20914 55022 20916 55074
rect 20412 54516 20468 54526
rect 20188 54460 20412 54516
rect 20412 54422 20468 54460
rect 19852 54292 19908 54302
rect 19740 53844 19796 53854
rect 19740 53750 19796 53788
rect 19628 53666 19684 53676
rect 19852 53730 19908 54236
rect 20860 54068 20916 55022
rect 21196 55074 21364 55076
rect 21196 55022 21310 55074
rect 21362 55022 21364 55074
rect 21196 55020 21364 55022
rect 21196 54514 21252 55020
rect 21308 55010 21364 55020
rect 21644 55074 21700 55086
rect 21644 55022 21646 55074
rect 21698 55022 21700 55074
rect 21196 54462 21198 54514
rect 21250 54462 21252 54514
rect 21196 54404 21252 54462
rect 20860 54002 20916 54012
rect 20972 54348 21196 54404
rect 19852 53678 19854 53730
rect 19906 53678 19908 53730
rect 19852 53666 19908 53678
rect 20300 53732 20356 53742
rect 19404 53508 19460 53518
rect 19404 53506 19572 53508
rect 19404 53454 19406 53506
rect 19458 53454 19572 53506
rect 19404 53452 19572 53454
rect 19404 53442 19460 53452
rect 18844 51314 18900 51324
rect 19068 52948 19124 52958
rect 19068 52274 19124 52892
rect 19292 52946 19348 53116
rect 19516 53060 19572 53452
rect 19628 53506 19684 53518
rect 19628 53454 19630 53506
rect 19682 53454 19684 53506
rect 19628 53284 19684 53454
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19628 53218 19684 53228
rect 19628 53060 19684 53070
rect 19516 53058 19684 53060
rect 19516 53006 19630 53058
rect 19682 53006 19684 53058
rect 19516 53004 19684 53006
rect 19628 52994 19684 53004
rect 19292 52894 19294 52946
rect 19346 52894 19348 52946
rect 19292 52882 19348 52894
rect 19852 52836 19908 52846
rect 19068 52222 19070 52274
rect 19122 52222 19124 52274
rect 19068 51378 19124 52222
rect 19180 52722 19236 52734
rect 19180 52670 19182 52722
rect 19234 52670 19236 52722
rect 19180 52612 19236 52670
rect 19180 52164 19236 52556
rect 19740 52724 19796 52734
rect 19852 52724 19908 52780
rect 19740 52722 19908 52724
rect 19740 52670 19742 52722
rect 19794 52670 19908 52722
rect 19740 52668 19908 52670
rect 19964 52722 20020 52734
rect 19964 52670 19966 52722
rect 20018 52670 20020 52722
rect 19740 52500 19796 52668
rect 19964 52612 20020 52670
rect 19964 52546 20020 52556
rect 20076 52722 20132 52734
rect 20076 52670 20078 52722
rect 20130 52670 20132 52722
rect 19516 52444 19796 52500
rect 19180 52098 19236 52108
rect 19404 52276 19460 52286
rect 19404 52162 19460 52220
rect 19404 52110 19406 52162
rect 19458 52110 19460 52162
rect 19404 52098 19460 52110
rect 19516 51604 19572 52444
rect 19628 52276 19684 52286
rect 20076 52276 20132 52670
rect 19628 52274 20132 52276
rect 19628 52222 19630 52274
rect 19682 52222 20132 52274
rect 19628 52220 20132 52222
rect 19628 51828 19684 52220
rect 19628 51762 19684 51772
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19516 51548 19796 51604
rect 19068 51326 19070 51378
rect 19122 51326 19124 51378
rect 19068 51314 19124 51326
rect 19180 51490 19236 51502
rect 19180 51438 19182 51490
rect 19234 51438 19236 51490
rect 19180 51380 19236 51438
rect 18732 51266 18788 51278
rect 18732 51214 18734 51266
rect 18786 51214 18788 51266
rect 18732 51156 18788 51214
rect 19180 51156 19236 51324
rect 18732 51100 19236 51156
rect 19292 51268 19348 51278
rect 18732 51044 18788 51100
rect 18732 50978 18788 50988
rect 18508 50764 19012 50820
rect 18396 49922 18452 50764
rect 18844 50596 18900 50606
rect 18956 50596 19012 50764
rect 18844 50594 19012 50596
rect 18844 50542 18846 50594
rect 18898 50542 19012 50594
rect 18844 50540 19012 50542
rect 18844 50530 18900 50540
rect 18396 49870 18398 49922
rect 18450 49870 18452 49922
rect 18396 49858 18452 49870
rect 18620 50482 18676 50494
rect 18620 50430 18622 50482
rect 18674 50430 18676 50482
rect 18620 49924 18676 50430
rect 18956 50370 19012 50382
rect 18956 50318 18958 50370
rect 19010 50318 19012 50370
rect 18956 50148 19012 50318
rect 18956 50082 19012 50092
rect 19180 50370 19236 50382
rect 19180 50318 19182 50370
rect 19234 50318 19236 50370
rect 18620 49858 18676 49868
rect 18956 49810 19012 49822
rect 18956 49758 18958 49810
rect 19010 49758 19012 49810
rect 18956 49700 19012 49758
rect 18956 49634 19012 49644
rect 18396 49140 18452 49150
rect 18284 49084 18396 49140
rect 18396 49074 18452 49084
rect 19068 49140 19124 49150
rect 18956 49028 19012 49038
rect 18508 48132 18564 48142
rect 18508 48038 18564 48076
rect 17724 47964 18116 48020
rect 17612 47572 17668 47582
rect 17388 47570 17668 47572
rect 17388 47518 17614 47570
rect 17666 47518 17668 47570
rect 17388 47516 17668 47518
rect 17276 47460 17332 47470
rect 17388 47460 17444 47516
rect 17612 47506 17668 47516
rect 17276 47458 17444 47460
rect 17276 47406 17278 47458
rect 17330 47406 17444 47458
rect 17276 47404 17444 47406
rect 17276 45668 17332 47404
rect 17724 47348 17780 47964
rect 17948 47796 18004 47806
rect 17612 47292 17780 47348
rect 17836 47348 17892 47358
rect 17500 47236 17556 47246
rect 17388 46452 17444 46462
rect 17388 46358 17444 46396
rect 17500 46228 17556 47180
rect 17388 46172 17556 46228
rect 17388 45890 17444 46172
rect 17388 45838 17390 45890
rect 17442 45838 17444 45890
rect 17388 45826 17444 45838
rect 17500 46004 17556 46014
rect 17500 45890 17556 45948
rect 17500 45838 17502 45890
rect 17554 45838 17556 45890
rect 17500 45826 17556 45838
rect 17612 45890 17668 47292
rect 17836 46900 17892 47292
rect 17948 47012 18004 47740
rect 18844 47796 18900 47806
rect 18956 47796 19012 48972
rect 19068 48804 19124 49084
rect 19180 48916 19236 50318
rect 19292 50034 19348 51212
rect 19628 51044 19684 51054
rect 19516 50818 19572 50830
rect 19516 50766 19518 50818
rect 19570 50766 19572 50818
rect 19516 50708 19572 50766
rect 19516 50642 19572 50652
rect 19628 50820 19684 50988
rect 19292 49982 19294 50034
rect 19346 49982 19348 50034
rect 19292 49970 19348 49982
rect 19404 50482 19460 50494
rect 19404 50430 19406 50482
rect 19458 50430 19460 50482
rect 19404 50036 19460 50430
rect 19516 50484 19572 50494
rect 19628 50484 19684 50764
rect 19516 50482 19684 50484
rect 19516 50430 19518 50482
rect 19570 50430 19684 50482
rect 19516 50428 19684 50430
rect 19516 50418 19572 50428
rect 19740 50372 19796 51548
rect 20188 51156 20244 51166
rect 20188 50706 20244 51100
rect 20188 50654 20190 50706
rect 20242 50654 20244 50706
rect 20188 50642 20244 50654
rect 19404 49970 19460 49980
rect 19628 50316 19796 50372
rect 20300 50372 20356 53676
rect 20412 53508 20468 53518
rect 20748 53508 20804 53518
rect 20468 53452 20692 53508
rect 20412 53414 20468 53452
rect 20524 53284 20580 53294
rect 20412 53228 20524 53284
rect 20636 53284 20692 53452
rect 20748 53414 20804 53452
rect 20636 53228 20804 53284
rect 20412 53170 20468 53228
rect 20524 53218 20580 53228
rect 20412 53118 20414 53170
rect 20466 53118 20468 53170
rect 20412 53106 20468 53118
rect 20636 53060 20692 53070
rect 20524 53058 20692 53060
rect 20524 53006 20638 53058
rect 20690 53006 20692 53058
rect 20524 53004 20692 53006
rect 20524 52500 20580 53004
rect 20636 52994 20692 53004
rect 20748 53058 20804 53228
rect 20748 53006 20750 53058
rect 20802 53006 20804 53058
rect 20748 52994 20804 53006
rect 20524 52434 20580 52444
rect 20636 52388 20692 52398
rect 20524 52052 20580 52062
rect 20524 51958 20580 51996
rect 20636 52050 20692 52332
rect 20860 52164 20916 52174
rect 20860 52070 20916 52108
rect 20636 51998 20638 52050
rect 20690 51998 20692 52050
rect 20636 51986 20692 51998
rect 20972 51380 21028 54348
rect 21196 54338 21252 54348
rect 21308 54626 21364 54638
rect 21308 54574 21310 54626
rect 21362 54574 21364 54626
rect 21308 54292 21364 54574
rect 21644 54628 21700 55022
rect 22204 55074 22260 55086
rect 22428 55076 22484 55086
rect 22204 55022 22206 55074
rect 22258 55022 22260 55074
rect 22204 54852 22260 55022
rect 22204 54786 22260 54796
rect 22316 55074 22484 55076
rect 22316 55022 22430 55074
rect 22482 55022 22484 55074
rect 22316 55020 22484 55022
rect 21644 54562 21700 54572
rect 21308 54226 21364 54236
rect 21420 54516 21476 54526
rect 21420 53842 21476 54460
rect 22204 54516 22260 54526
rect 22316 54516 22372 55020
rect 22428 55010 22484 55020
rect 22764 55076 22820 55086
rect 23324 55076 23380 55086
rect 22764 55074 22932 55076
rect 22764 55022 22766 55074
rect 22818 55022 22932 55074
rect 22764 55020 22932 55022
rect 22764 55010 22820 55020
rect 22764 54852 22820 54862
rect 22260 54460 22372 54516
rect 22428 54628 22484 54638
rect 22428 54514 22484 54572
rect 22428 54462 22430 54514
rect 22482 54462 22484 54514
rect 22204 54422 22260 54460
rect 22428 54450 22484 54462
rect 21420 53790 21422 53842
rect 21474 53790 21476 53842
rect 21420 53778 21476 53790
rect 21532 54404 21588 54414
rect 21196 52836 21252 52846
rect 21196 52742 21252 52780
rect 21420 52388 21476 52398
rect 20636 51378 21028 51380
rect 20636 51326 20974 51378
rect 21026 51326 21028 51378
rect 20636 51324 21028 51326
rect 19628 49924 19684 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19628 49830 19684 49868
rect 19404 49810 19460 49822
rect 19404 49758 19406 49810
rect 19458 49758 19460 49810
rect 19292 49252 19348 49262
rect 19292 49138 19348 49196
rect 19292 49086 19294 49138
rect 19346 49086 19348 49138
rect 19292 49074 19348 49086
rect 19292 48916 19348 48926
rect 19180 48860 19292 48916
rect 19292 48850 19348 48860
rect 19068 48748 19236 48804
rect 18900 47740 19012 47796
rect 18844 47730 18900 47740
rect 18732 47460 18788 47470
rect 18732 47458 18900 47460
rect 18732 47406 18734 47458
rect 18786 47406 18900 47458
rect 18732 47404 18900 47406
rect 18732 47394 18788 47404
rect 18508 47348 18564 47358
rect 18396 47346 18564 47348
rect 18396 47294 18510 47346
rect 18562 47294 18564 47346
rect 18396 47292 18564 47294
rect 18172 47236 18228 47246
rect 18396 47236 18452 47292
rect 18508 47282 18564 47292
rect 18172 47234 18340 47236
rect 18172 47182 18174 47234
rect 18226 47182 18340 47234
rect 18172 47180 18340 47182
rect 18172 47170 18228 47180
rect 18004 46956 18228 47012
rect 17948 46946 18004 46956
rect 17724 46844 17892 46900
rect 17724 46674 17780 46844
rect 18060 46788 18116 46798
rect 18060 46694 18116 46732
rect 17724 46622 17726 46674
rect 17778 46622 17780 46674
rect 17724 46564 17780 46622
rect 17836 46676 17892 46686
rect 17836 46582 17892 46620
rect 17724 46116 17780 46508
rect 17948 46562 18004 46574
rect 17948 46510 17950 46562
rect 18002 46510 18004 46562
rect 17948 46116 18004 46510
rect 17724 46060 17892 46116
rect 17612 45838 17614 45890
rect 17666 45838 17668 45890
rect 17612 45826 17668 45838
rect 17724 45892 17780 45902
rect 17724 45798 17780 45836
rect 17276 45612 17668 45668
rect 17388 45444 17444 45454
rect 17388 45332 17444 45388
rect 17388 45330 17556 45332
rect 17388 45278 17390 45330
rect 17442 45278 17556 45330
rect 17388 45276 17556 45278
rect 17388 45266 17444 45276
rect 16828 43652 17220 43708
rect 17388 44548 17444 44558
rect 16828 43650 16884 43652
rect 16828 43598 16830 43650
rect 16882 43598 16884 43650
rect 16828 43586 16884 43598
rect 16940 43540 16996 43550
rect 16604 42866 16772 42868
rect 16604 42814 16606 42866
rect 16658 42814 16772 42866
rect 16604 42812 16772 42814
rect 16828 42868 16884 42878
rect 16604 42644 16660 42812
rect 16604 42578 16660 42588
rect 16828 42082 16884 42812
rect 16828 42030 16830 42082
rect 16882 42030 16884 42082
rect 16604 41972 16660 41982
rect 16604 41970 16772 41972
rect 16604 41918 16606 41970
rect 16658 41918 16772 41970
rect 16604 41916 16772 41918
rect 16604 41906 16660 41916
rect 16716 40740 16772 41916
rect 16828 41186 16884 42030
rect 16828 41134 16830 41186
rect 16882 41134 16884 41186
rect 16828 41122 16884 41134
rect 16716 40626 16772 40684
rect 16716 40574 16718 40626
rect 16770 40574 16772 40626
rect 16716 40562 16772 40574
rect 16492 40516 16548 40526
rect 16492 40422 16548 40460
rect 16828 40402 16884 40414
rect 16828 40350 16830 40402
rect 16882 40350 16884 40402
rect 16380 40236 16660 40292
rect 16380 39620 16436 39630
rect 16380 39618 16548 39620
rect 16380 39566 16382 39618
rect 16434 39566 16548 39618
rect 16380 39564 16548 39566
rect 16380 39554 16436 39564
rect 16156 39340 16436 39396
rect 16044 39228 16324 39284
rect 16156 39060 16212 39070
rect 15708 38834 15764 38846
rect 15708 38782 15710 38834
rect 15762 38782 15764 38834
rect 15708 38164 15764 38782
rect 16044 38836 16100 38846
rect 16044 38722 16100 38780
rect 16156 38834 16212 39004
rect 16156 38782 16158 38834
rect 16210 38782 16212 38834
rect 16156 38770 16212 38782
rect 16044 38670 16046 38722
rect 16098 38670 16100 38722
rect 15932 38276 15988 38286
rect 15932 38182 15988 38220
rect 15708 35810 15764 38108
rect 16044 38052 16100 38670
rect 16044 37986 16100 37996
rect 15820 37492 15876 37502
rect 15820 37268 15876 37436
rect 15820 37202 15876 37212
rect 16044 37268 16100 37278
rect 16044 37174 16100 37212
rect 15820 36484 15876 36494
rect 15820 36390 15876 36428
rect 15708 35758 15710 35810
rect 15762 35758 15764 35810
rect 15708 35746 15764 35758
rect 15372 34974 15374 35026
rect 15426 34974 15428 35026
rect 15372 34962 15428 34974
rect 16044 35698 16100 35710
rect 16044 35646 16046 35698
rect 16098 35646 16100 35698
rect 16044 34916 16100 35646
rect 16044 34822 16100 34860
rect 15708 34356 15764 34366
rect 15260 34300 15540 34356
rect 15148 34020 15204 34030
rect 15148 34018 15316 34020
rect 15148 33966 15150 34018
rect 15202 33966 15316 34018
rect 15148 33964 15316 33966
rect 15148 33954 15204 33964
rect 14812 33406 14814 33458
rect 14866 33406 14868 33458
rect 14812 33394 14868 33406
rect 14700 33170 14756 33180
rect 15148 32676 15204 32686
rect 15260 32676 15316 33964
rect 15372 33908 15428 33918
rect 15372 33814 15428 33852
rect 15372 32900 15428 32910
rect 15484 32900 15540 34300
rect 15708 34262 15764 34300
rect 16268 34130 16324 39228
rect 16268 34078 16270 34130
rect 16322 34078 16324 34130
rect 16268 34066 16324 34078
rect 15596 33236 15652 33246
rect 15596 33142 15652 33180
rect 15428 32844 15540 32900
rect 15372 32834 15428 32844
rect 15932 32788 15988 32798
rect 15932 32694 15988 32732
rect 14588 32498 14644 32508
rect 14812 32620 15148 32676
rect 15204 32620 15316 32676
rect 15708 32676 15764 32686
rect 14812 32562 14868 32620
rect 15148 32582 15204 32620
rect 15708 32582 15764 32620
rect 14812 32510 14814 32562
rect 14866 32510 14868 32562
rect 14812 32498 14868 32510
rect 15596 32562 15652 32574
rect 15596 32510 15598 32562
rect 15650 32510 15652 32562
rect 15148 32452 15204 32462
rect 15148 32358 15204 32396
rect 14700 31892 14756 31902
rect 14700 31798 14756 31836
rect 14364 31490 14420 31500
rect 14700 31668 14756 31678
rect 14476 31220 14532 31230
rect 14252 31218 14532 31220
rect 14252 31166 14478 31218
rect 14530 31166 14532 31218
rect 14252 31164 14532 31166
rect 14476 31154 14532 31164
rect 8540 31042 8596 31052
rect 9548 31108 9604 31118
rect 9100 30436 9156 30446
rect 9100 30210 9156 30380
rect 9100 30158 9102 30210
rect 9154 30158 9156 30210
rect 9100 30146 9156 30158
rect 9548 29988 9604 31052
rect 9772 30994 9828 31006
rect 9772 30942 9774 30994
rect 9826 30942 9828 30994
rect 9660 29988 9716 29998
rect 9548 29986 9716 29988
rect 9548 29934 9662 29986
rect 9714 29934 9716 29986
rect 9548 29932 9716 29934
rect 9660 29922 9716 29932
rect 8316 29586 8372 29596
rect 5628 28530 6020 28532
rect 5628 28478 5966 28530
rect 6018 28478 6020 28530
rect 5628 28476 6020 28478
rect 1708 28420 1764 28430
rect 1708 28326 1764 28364
rect 2044 28084 2100 28094
rect 2044 27990 2100 28028
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27636 1764 27806
rect 5628 27858 5684 28476
rect 5964 28466 6020 28476
rect 6300 28642 6356 28654
rect 6300 28590 6302 28642
rect 6354 28590 6356 28642
rect 5628 27806 5630 27858
rect 5682 27806 5684 27858
rect 5628 27794 5684 27806
rect 6076 27860 6132 27870
rect 6076 27766 6132 27804
rect 1708 27570 1764 27580
rect 2492 27746 2548 27758
rect 2492 27694 2494 27746
rect 2546 27694 2548 27746
rect 2492 27636 2548 27694
rect 2492 27570 2548 27580
rect 2044 27524 2100 27534
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1708 26964 1764 26974
rect 1708 26402 1764 26908
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 26338 1764 26350
rect 1932 26292 1988 27134
rect 2044 26514 2100 27468
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27074 4340 27086
rect 4284 27022 4286 27074
rect 4338 27022 4340 27074
rect 2044 26462 2046 26514
rect 2098 26462 2100 26514
rect 2044 26450 2100 26462
rect 2492 26964 2548 26974
rect 2268 26292 2324 26302
rect 1932 26226 1988 26236
rect 2044 26236 2268 26292
rect 1708 25394 1764 25406
rect 1708 25342 1710 25394
rect 1762 25342 1764 25394
rect 1708 24948 1764 25342
rect 2044 25394 2100 26236
rect 2268 26226 2324 26236
rect 2380 26290 2436 26302
rect 2380 26238 2382 26290
rect 2434 26238 2436 26290
rect 2380 26180 2436 26238
rect 2380 25620 2436 26124
rect 2380 25554 2436 25564
rect 2492 25618 2548 26908
rect 2716 26516 2772 26526
rect 2716 26422 2772 26460
rect 3164 26180 3220 26190
rect 3164 26086 3220 26124
rect 4284 26068 4340 27022
rect 6300 26852 6356 28590
rect 8316 27972 8372 27982
rect 5068 26628 5124 26638
rect 5068 26514 5124 26572
rect 5068 26462 5070 26514
rect 5122 26462 5124 26514
rect 4396 26292 4452 26302
rect 4396 26198 4452 26236
rect 4844 26292 4900 26302
rect 4844 26198 4900 26236
rect 4284 26002 4340 26012
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 2492 25566 2494 25618
rect 2546 25566 2548 25618
rect 2492 25554 2548 25566
rect 2044 25342 2046 25394
rect 2098 25342 2100 25394
rect 2044 25330 2100 25342
rect 4172 25506 4228 25518
rect 4172 25454 4174 25506
rect 4226 25454 4228 25506
rect 1708 24882 1764 24892
rect 2940 25282 2996 25294
rect 2940 25230 2942 25282
rect 2994 25230 2996 25282
rect 2940 24948 2996 25230
rect 4172 25284 4228 25454
rect 5068 25506 5124 26462
rect 5740 26628 5796 26638
rect 5516 26290 5572 26302
rect 5516 26238 5518 26290
rect 5570 26238 5572 26290
rect 5516 25732 5572 26238
rect 5068 25454 5070 25506
rect 5122 25454 5124 25506
rect 5068 25442 5124 25454
rect 5180 25676 5516 25732
rect 4396 25396 4452 25406
rect 4396 25302 4452 25340
rect 5180 25396 5236 25676
rect 5516 25666 5572 25676
rect 5740 25618 5796 26572
rect 5964 26292 6020 26302
rect 5964 26290 6244 26292
rect 5964 26238 5966 26290
rect 6018 26238 6244 26290
rect 5964 26236 6244 26238
rect 5964 26226 6020 26236
rect 5740 25566 5742 25618
rect 5794 25566 5796 25618
rect 5740 25554 5796 25566
rect 4172 25218 4228 25228
rect 4732 25284 4788 25294
rect 4732 25190 4788 25228
rect 2940 24882 2996 24892
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 5068 24724 5124 24734
rect 5180 24724 5236 25340
rect 6188 25394 6244 26236
rect 6188 25342 6190 25394
rect 6242 25342 6244 25394
rect 6188 25330 6244 25342
rect 6300 25284 6356 26796
rect 8204 27970 8372 27972
rect 8204 27918 8318 27970
rect 8370 27918 8372 27970
rect 8204 27916 8372 27918
rect 8204 26402 8260 27916
rect 8316 27906 8372 27916
rect 9548 27860 9604 27870
rect 9436 27858 9604 27860
rect 9436 27806 9550 27858
rect 9602 27806 9604 27858
rect 9436 27804 9604 27806
rect 9100 27636 9156 27646
rect 8988 27634 9156 27636
rect 8988 27582 9102 27634
rect 9154 27582 9156 27634
rect 8988 27580 9156 27582
rect 8876 27188 8932 27198
rect 8876 27074 8932 27132
rect 8876 27022 8878 27074
rect 8930 27022 8932 27074
rect 8876 27010 8932 27022
rect 8988 26908 9044 27580
rect 9100 27570 9156 27580
rect 8204 26350 8206 26402
rect 8258 26350 8260 26402
rect 8204 26180 8260 26350
rect 6524 25620 6580 25630
rect 6524 25506 6580 25564
rect 6524 25454 6526 25506
rect 6578 25454 6580 25506
rect 6524 25442 6580 25454
rect 6300 25218 6356 25228
rect 5964 25172 6020 25182
rect 5068 24722 5236 24724
rect 5068 24670 5070 24722
rect 5122 24670 5236 24722
rect 5068 24668 5236 24670
rect 5516 24722 5572 24734
rect 5516 24670 5518 24722
rect 5570 24670 5572 24722
rect 5068 24658 5124 24668
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 5516 23828 5572 24670
rect 5964 23938 6020 25116
rect 7756 24724 7812 24734
rect 8204 24724 8260 26124
rect 8876 26852 9044 26908
rect 9212 27412 9268 27422
rect 9212 26962 9268 27356
rect 9212 26910 9214 26962
rect 9266 26910 9268 26962
rect 9212 26898 9268 26910
rect 8764 25732 8820 25742
rect 8764 25506 8820 25676
rect 8764 25454 8766 25506
rect 8818 25454 8820 25506
rect 8764 25442 8820 25454
rect 7756 24722 8260 24724
rect 7756 24670 7758 24722
rect 7810 24670 8260 24722
rect 7756 24668 8260 24670
rect 7756 24658 7812 24668
rect 5964 23886 5966 23938
rect 6018 23886 6020 23938
rect 5964 23874 6020 23886
rect 7980 24500 8036 24510
rect 5628 23828 5684 23838
rect 5516 23826 5684 23828
rect 5516 23774 5630 23826
rect 5682 23774 5684 23826
rect 5516 23772 5684 23774
rect 5628 23762 5684 23772
rect 1932 23538 1988 23548
rect 7308 23716 7364 23726
rect 4172 23380 4228 23390
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22484 1988 22494
rect 1932 22390 1988 22428
rect 4172 22370 4228 23324
rect 4284 23268 4340 23278
rect 4284 23154 4340 23212
rect 4284 23102 4286 23154
rect 4338 23102 4340 23154
rect 4284 23090 4340 23102
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 22318 4174 22370
rect 4226 22318 4228 22370
rect 4172 22306 4228 22318
rect 6300 22260 6356 22270
rect 4284 21812 4340 21822
rect 4284 21586 4340 21756
rect 6300 21812 6356 22204
rect 6860 22148 6916 22158
rect 6748 21812 6804 21822
rect 6300 21810 6580 21812
rect 6300 21758 6302 21810
rect 6354 21758 6580 21810
rect 6300 21756 6580 21758
rect 6300 21746 6356 21756
rect 4284 21534 4286 21586
rect 4338 21534 4340 21586
rect 4284 21522 4340 21534
rect 5964 21588 6020 21598
rect 1932 21476 1988 21486
rect 1932 21382 1988 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5852 20804 5908 20814
rect 5852 20710 5908 20748
rect 3276 20468 3332 20478
rect 1708 19012 1764 19022
rect 1708 18918 1764 18956
rect 1708 17442 1764 17454
rect 1708 17390 1710 17442
rect 1762 17390 1764 17442
rect 1708 16884 1764 17390
rect 1708 16818 1764 16828
rect 3276 9604 3332 20412
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 5964 19234 6020 21532
rect 6076 20580 6132 20590
rect 6412 20580 6468 20590
rect 6076 20578 6468 20580
rect 6076 20526 6078 20578
rect 6130 20526 6414 20578
rect 6466 20526 6468 20578
rect 6076 20524 6468 20526
rect 6076 20514 6132 20524
rect 6300 20356 6356 20366
rect 6076 19908 6132 19918
rect 6076 19814 6132 19852
rect 5964 19182 5966 19234
rect 6018 19182 6020 19234
rect 5964 19124 6020 19182
rect 5964 19068 6244 19124
rect 5740 18564 5796 18574
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5404 17108 5460 17118
rect 5404 17014 5460 17052
rect 5740 16770 5796 18508
rect 5740 16718 5742 16770
rect 5794 16718 5796 16770
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5740 15988 5796 16718
rect 6076 16994 6132 17006
rect 6076 16942 6078 16994
rect 6130 16942 6132 16994
rect 6076 16884 6132 16942
rect 5852 16548 5908 16558
rect 5852 16210 5908 16492
rect 5852 16158 5854 16210
rect 5906 16158 5908 16210
rect 5852 16146 5908 16158
rect 5740 15922 5796 15932
rect 6076 15874 6132 16828
rect 6076 15822 6078 15874
rect 6130 15822 6132 15874
rect 6076 15764 6132 15822
rect 5852 15708 6132 15764
rect 5628 15316 5684 15326
rect 5628 15222 5684 15260
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 5852 12180 5908 15708
rect 6188 15652 6244 19068
rect 5964 15596 6244 15652
rect 5964 13970 6020 15596
rect 5964 13918 5966 13970
rect 6018 13918 6020 13970
rect 5964 13524 6020 13918
rect 5964 13458 6020 13468
rect 6076 15202 6132 15214
rect 6076 15150 6078 15202
rect 6130 15150 6132 15202
rect 5740 12178 5908 12180
rect 5740 12126 5854 12178
rect 5906 12126 5908 12178
rect 5740 12124 5908 12126
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5740 10610 5796 12124
rect 5852 12114 5908 12124
rect 6076 10724 6132 15150
rect 6300 14756 6356 20300
rect 6412 20020 6468 20524
rect 6412 19234 6468 19964
rect 6412 19182 6414 19234
rect 6466 19182 6468 19234
rect 6412 19170 6468 19182
rect 6524 18452 6580 21756
rect 6748 21586 6804 21756
rect 6748 21534 6750 21586
rect 6802 21534 6804 21586
rect 6748 21522 6804 21534
rect 6748 20580 6804 20590
rect 6860 20580 6916 22092
rect 6972 21698 7028 21710
rect 6972 21646 6974 21698
rect 7026 21646 7028 21698
rect 6972 21588 7028 21646
rect 6972 21522 7028 21532
rect 6748 20578 6916 20580
rect 6748 20526 6750 20578
rect 6802 20526 6916 20578
rect 6748 20524 6916 20526
rect 6748 20514 6804 20524
rect 6748 19908 6804 19918
rect 6748 18564 6804 19852
rect 6748 18470 6804 18508
rect 6412 16996 6468 17006
rect 6412 16098 6468 16940
rect 6524 16994 6580 18396
rect 6524 16942 6526 16994
rect 6578 16942 6580 16994
rect 6524 16930 6580 16942
rect 6412 16046 6414 16098
rect 6466 16046 6468 16098
rect 6412 16034 6468 16046
rect 6524 15988 6580 15998
rect 6524 15314 6580 15932
rect 6524 15262 6526 15314
rect 6578 15262 6580 15314
rect 6524 15250 6580 15262
rect 6748 15874 6804 15886
rect 6748 15822 6750 15874
rect 6802 15822 6804 15874
rect 6300 14690 6356 14700
rect 6636 15202 6692 15214
rect 6636 15150 6638 15202
rect 6690 15150 6692 15202
rect 6188 14532 6244 14542
rect 6188 14438 6244 14476
rect 6636 14530 6692 15150
rect 6748 14644 6804 15822
rect 6860 15148 6916 20524
rect 7084 20580 7140 20590
rect 7084 20578 7252 20580
rect 7084 20526 7086 20578
rect 7138 20526 7252 20578
rect 7084 20524 7252 20526
rect 7084 20514 7140 20524
rect 7084 20020 7140 20030
rect 7084 19926 7140 19964
rect 7196 19796 7252 20524
rect 7308 20018 7364 23660
rect 7868 23268 7924 23278
rect 7868 23154 7924 23212
rect 7868 23102 7870 23154
rect 7922 23102 7924 23154
rect 7420 21812 7476 21822
rect 7420 20802 7476 21756
rect 7420 20750 7422 20802
rect 7474 20750 7476 20802
rect 7420 20738 7476 20750
rect 7868 20804 7924 23102
rect 7980 23042 8036 24444
rect 8764 24500 8820 24510
rect 8764 24406 8820 24444
rect 8764 23380 8820 23390
rect 8316 23156 8372 23166
rect 8764 23156 8820 23324
rect 8876 23268 8932 26852
rect 9436 26740 9492 27804
rect 9548 27794 9604 27804
rect 9660 27412 9716 27422
rect 9660 27074 9716 27356
rect 9660 27022 9662 27074
rect 9714 27022 9716 27074
rect 9660 27010 9716 27022
rect 9772 26964 9828 30942
rect 12572 30996 12628 31006
rect 13020 30996 13076 31006
rect 12572 30994 13076 30996
rect 12572 30942 12574 30994
rect 12626 30942 13022 30994
rect 13074 30942 13076 30994
rect 12572 30940 13076 30942
rect 12572 30436 12628 30940
rect 13020 30930 13076 30940
rect 12572 30370 12628 30380
rect 14588 30436 14644 30446
rect 12236 30212 12292 30222
rect 12572 30212 12628 30222
rect 12236 30118 12292 30156
rect 12460 30210 12628 30212
rect 12460 30158 12574 30210
rect 12626 30158 12628 30210
rect 12460 30156 12628 30158
rect 11788 29652 11844 29662
rect 11788 29558 11844 29596
rect 12348 29652 12404 29662
rect 10108 29428 10164 29438
rect 10108 28196 10164 29372
rect 12348 29426 12404 29596
rect 12348 29374 12350 29426
rect 12402 29374 12404 29426
rect 12348 29362 12404 29374
rect 9884 28140 10388 28196
rect 9884 28082 9940 28140
rect 9884 28030 9886 28082
rect 9938 28030 9940 28082
rect 9884 28018 9940 28030
rect 10332 27188 10388 28140
rect 12460 27188 12516 30156
rect 12572 30146 12628 30156
rect 12572 29316 12628 29326
rect 13020 29316 13076 29326
rect 12572 29222 12628 29260
rect 12684 29314 13076 29316
rect 12684 29262 13022 29314
rect 13074 29262 13076 29314
rect 12684 29260 13076 29262
rect 12684 28642 12740 29260
rect 13020 29250 13076 29260
rect 12684 28590 12686 28642
rect 12738 28590 12740 28642
rect 12684 28578 12740 28590
rect 12908 28644 12964 28654
rect 12908 28530 12964 28588
rect 12908 28478 12910 28530
rect 12962 28478 12964 28530
rect 12908 28466 12964 28478
rect 13468 28642 13524 28654
rect 13468 28590 13470 28642
rect 13522 28590 13524 28642
rect 10332 27094 10388 27132
rect 12348 27132 12516 27188
rect 9884 26964 9940 26974
rect 9772 26962 10052 26964
rect 9772 26910 9886 26962
rect 9938 26910 10052 26962
rect 9772 26908 10052 26910
rect 9884 26898 9940 26908
rect 9996 26852 10500 26908
rect 12124 26852 12180 26862
rect 9436 26674 9492 26684
rect 10444 26516 10500 26852
rect 11788 26850 12180 26852
rect 11788 26798 12126 26850
rect 12178 26798 12180 26850
rect 11788 26796 12180 26798
rect 11340 26740 11396 26750
rect 9660 26404 9716 26414
rect 9212 26402 9716 26404
rect 9212 26350 9662 26402
rect 9714 26350 9716 26402
rect 9212 26348 9716 26350
rect 8988 26066 9044 26078
rect 8988 26014 8990 26066
rect 9042 26014 9044 26066
rect 8988 23716 9044 26014
rect 9212 25506 9268 26348
rect 9660 26338 9716 26348
rect 9996 26404 10052 26414
rect 9996 26310 10052 26348
rect 10444 26290 10500 26460
rect 10444 26238 10446 26290
rect 10498 26238 10500 26290
rect 10444 26226 10500 26238
rect 11228 26684 11340 26740
rect 11228 26290 11284 26684
rect 11340 26674 11396 26684
rect 11228 26238 11230 26290
rect 11282 26238 11284 26290
rect 11228 26226 11284 26238
rect 11788 26290 11844 26796
rect 12124 26786 12180 26796
rect 11788 26238 11790 26290
rect 11842 26238 11844 26290
rect 11788 26226 11844 26238
rect 10780 26180 10836 26190
rect 10780 26086 10836 26124
rect 11340 26180 11396 26190
rect 9212 25454 9214 25506
rect 9266 25454 9268 25506
rect 9212 25442 9268 25454
rect 11340 25506 11396 26124
rect 12348 25732 12404 27132
rect 12460 26964 12516 26974
rect 12460 26870 12516 26908
rect 13468 26740 13524 28590
rect 13916 28644 13972 28654
rect 13916 28550 13972 28588
rect 14588 26908 14644 30380
rect 14700 29988 14756 31612
rect 15596 31668 15652 32510
rect 14812 30994 14868 31006
rect 14812 30942 14814 30994
rect 14866 30942 14868 30994
rect 14812 30212 14868 30942
rect 15596 30884 15652 31612
rect 16380 31332 16436 39340
rect 16492 38948 16548 39564
rect 16604 39396 16660 40236
rect 16828 40180 16884 40350
rect 16828 40068 16884 40124
rect 16716 40012 16884 40068
rect 16716 39620 16772 40012
rect 16828 39844 16884 39854
rect 16828 39750 16884 39788
rect 16716 39564 16884 39620
rect 16604 39340 16772 39396
rect 16604 38948 16660 38958
rect 16492 38892 16604 38948
rect 16604 38882 16660 38892
rect 16716 38946 16772 39340
rect 16828 39284 16884 39564
rect 16828 39218 16884 39228
rect 16716 38894 16718 38946
rect 16770 38894 16772 38946
rect 16716 38882 16772 38894
rect 16492 38052 16548 38062
rect 16492 36482 16548 37996
rect 16604 37940 16660 37950
rect 16604 37938 16772 37940
rect 16604 37886 16606 37938
rect 16658 37886 16772 37938
rect 16604 37884 16772 37886
rect 16604 37874 16660 37884
rect 16492 36430 16494 36482
rect 16546 36430 16548 36482
rect 16492 36418 16548 36430
rect 16716 36484 16772 37884
rect 16716 36390 16772 36428
rect 16828 37156 16884 37166
rect 16940 37156 16996 43484
rect 16828 37154 16996 37156
rect 16828 37102 16830 37154
rect 16882 37102 16996 37154
rect 16828 37100 16996 37102
rect 17052 42644 17108 43652
rect 17388 43428 17444 44492
rect 17500 44212 17556 45276
rect 17500 44146 17556 44156
rect 17612 44660 17668 45612
rect 17836 45388 17892 46060
rect 17948 46050 18004 46060
rect 17948 45892 18004 45902
rect 17948 45798 18004 45836
rect 17836 45332 18004 45388
rect 17612 43988 17668 44604
rect 17724 45108 17780 45118
rect 17724 44100 17780 45052
rect 17836 44994 17892 45006
rect 17836 44942 17838 44994
rect 17890 44942 17892 44994
rect 17836 44324 17892 44942
rect 17836 44258 17892 44268
rect 17724 44034 17780 44044
rect 17948 44100 18004 45332
rect 18172 45220 18228 46956
rect 18284 46228 18340 47180
rect 18396 47170 18452 47180
rect 18620 47236 18676 47246
rect 18508 47124 18564 47134
rect 18508 47012 18564 47068
rect 18508 46676 18564 46956
rect 18508 46610 18564 46620
rect 18284 46162 18340 46172
rect 18508 46116 18564 46126
rect 18284 46004 18340 46014
rect 18284 45332 18340 45948
rect 18508 45778 18564 46060
rect 18620 46114 18676 47180
rect 18844 47068 18900 47404
rect 18732 47012 18900 47068
rect 19068 47458 19124 47470
rect 19068 47406 19070 47458
rect 19122 47406 19124 47458
rect 19068 47124 19124 47406
rect 18732 46564 18788 47012
rect 19068 46898 19124 47068
rect 19068 46846 19070 46898
rect 19122 46846 19124 46898
rect 19068 46834 19124 46846
rect 18844 46788 18900 46798
rect 18844 46786 19012 46788
rect 18844 46734 18846 46786
rect 18898 46734 19012 46786
rect 18844 46732 19012 46734
rect 18844 46722 18900 46732
rect 18732 46508 18900 46564
rect 18620 46062 18622 46114
rect 18674 46062 18676 46114
rect 18620 45892 18676 46062
rect 18620 45826 18676 45836
rect 18732 46228 18788 46238
rect 18508 45726 18510 45778
rect 18562 45726 18564 45778
rect 18508 45714 18564 45726
rect 18396 45332 18452 45342
rect 18340 45330 18452 45332
rect 18340 45278 18398 45330
rect 18450 45278 18452 45330
rect 18340 45276 18452 45278
rect 18284 45238 18340 45276
rect 18396 45266 18452 45276
rect 17948 44034 18004 44044
rect 18060 45164 18228 45220
rect 17276 43372 17444 43428
rect 17500 43932 17668 43988
rect 17500 43650 17556 43932
rect 17500 43598 17502 43650
rect 17554 43598 17556 43650
rect 17500 43428 17556 43598
rect 17612 43652 17668 43662
rect 17612 43558 17668 43596
rect 17724 43540 17780 43550
rect 17724 43446 17780 43484
rect 17500 43372 17668 43428
rect 17164 42644 17220 42654
rect 17052 42642 17220 42644
rect 17052 42590 17166 42642
rect 17218 42590 17220 42642
rect 17052 42588 17220 42590
rect 16604 35588 16660 35598
rect 16828 35588 16884 37100
rect 16604 35586 16884 35588
rect 16604 35534 16606 35586
rect 16658 35534 16884 35586
rect 16604 35532 16884 35534
rect 16604 35476 16660 35532
rect 16604 35410 16660 35420
rect 16492 34804 16548 34814
rect 16492 34244 16548 34748
rect 16828 34692 16884 34702
rect 16828 34354 16884 34636
rect 16828 34302 16830 34354
rect 16882 34302 16884 34354
rect 16828 34290 16884 34302
rect 16492 34178 16548 34188
rect 17052 33572 17108 42588
rect 17164 42578 17220 42588
rect 17276 42420 17332 43372
rect 17388 42978 17444 42990
rect 17388 42926 17390 42978
rect 17442 42926 17444 42978
rect 17388 42868 17444 42926
rect 17388 42802 17444 42812
rect 17164 42364 17332 42420
rect 17388 42644 17444 42654
rect 17164 39844 17220 42364
rect 17388 41972 17444 42588
rect 17164 39778 17220 39788
rect 17276 41412 17332 41422
rect 17276 41188 17332 41356
rect 17276 39620 17332 41132
rect 17164 39618 17332 39620
rect 17164 39566 17278 39618
rect 17330 39566 17332 39618
rect 17164 39564 17332 39566
rect 17164 38052 17220 39564
rect 17276 39554 17332 39564
rect 17388 40290 17444 41916
rect 17388 40238 17390 40290
rect 17442 40238 17444 40290
rect 17388 39058 17444 40238
rect 17500 40404 17556 40414
rect 17500 40290 17556 40348
rect 17500 40238 17502 40290
rect 17554 40238 17556 40290
rect 17500 40226 17556 40238
rect 17612 39508 17668 43372
rect 18060 41972 18116 45164
rect 18172 44996 18228 45006
rect 18172 42868 18228 44940
rect 18732 43764 18788 46172
rect 18844 46116 18900 46508
rect 18844 46050 18900 46060
rect 18844 45892 18900 45902
rect 18844 45668 18900 45836
rect 18844 45602 18900 45612
rect 18956 45444 19012 46732
rect 19180 46676 19236 48748
rect 19292 48130 19348 48142
rect 19292 48078 19294 48130
rect 19346 48078 19348 48130
rect 19292 47460 19348 48078
rect 19292 47394 19348 47404
rect 19068 46620 19236 46676
rect 19404 47236 19460 49758
rect 20188 49810 20244 49822
rect 20188 49758 20190 49810
rect 20242 49758 20244 49810
rect 20188 49588 20244 49758
rect 20188 49522 20244 49532
rect 19740 49250 19796 49262
rect 19740 49198 19742 49250
rect 19794 49198 19796 49250
rect 19740 48804 19796 49198
rect 20300 49028 20356 50316
rect 20524 50482 20580 50494
rect 20524 50430 20526 50482
rect 20578 50430 20580 50482
rect 20300 48962 20356 48972
rect 20412 49922 20468 49934
rect 20412 49870 20414 49922
rect 20466 49870 20468 49922
rect 19740 48748 20244 48804
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48354 20244 48748
rect 20188 48302 20190 48354
rect 20242 48302 20244 48354
rect 20188 48290 20244 48302
rect 20412 48242 20468 49870
rect 20524 49588 20580 50430
rect 20636 50482 20692 51324
rect 20972 51314 21028 51324
rect 21308 52276 21364 52286
rect 20972 50820 21028 50830
rect 20636 50430 20638 50482
rect 20690 50430 20692 50482
rect 20636 50418 20692 50430
rect 20860 50484 20916 50522
rect 20860 50418 20916 50428
rect 20524 49522 20580 49532
rect 20748 49140 20804 49150
rect 20748 49046 20804 49084
rect 20412 48190 20414 48242
rect 20466 48190 20468 48242
rect 20188 48020 20244 48030
rect 19628 47572 19684 47610
rect 19628 47506 19684 47516
rect 19740 47348 19796 47358
rect 19740 47254 19796 47292
rect 19404 46674 19460 47180
rect 19516 47234 19572 47246
rect 19516 47182 19518 47234
rect 19570 47182 19572 47234
rect 19516 47012 19572 47182
rect 19516 46946 19572 46956
rect 19628 47124 19684 47134
rect 19628 46900 19684 47068
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19628 46834 19684 46844
rect 19404 46622 19406 46674
rect 19458 46622 19460 46674
rect 19068 45668 19124 46620
rect 19404 46610 19460 46622
rect 19852 46674 19908 46686
rect 19852 46622 19854 46674
rect 19906 46622 19908 46674
rect 19180 46452 19236 46462
rect 19852 46452 19908 46622
rect 19180 46450 19908 46452
rect 19180 46398 19182 46450
rect 19234 46398 19908 46450
rect 19180 46396 19908 46398
rect 19180 46386 19236 46396
rect 19964 46228 20020 46238
rect 19964 46114 20020 46172
rect 19964 46062 19966 46114
rect 20018 46062 20020 46114
rect 19964 46050 20020 46062
rect 19740 45892 19796 45902
rect 19292 45890 19796 45892
rect 19292 45838 19742 45890
rect 19794 45838 19796 45890
rect 19292 45836 19796 45838
rect 19292 45668 19348 45836
rect 19740 45826 19796 45836
rect 20076 45892 20132 45930
rect 20188 45892 20244 47964
rect 20300 47236 20356 47246
rect 20300 47142 20356 47180
rect 20300 46900 20356 46910
rect 20300 46562 20356 46844
rect 20300 46510 20302 46562
rect 20354 46510 20356 46562
rect 20300 46498 20356 46510
rect 20412 46452 20468 48190
rect 20748 48132 20804 48142
rect 20636 47460 20692 47470
rect 20524 47348 20580 47358
rect 20524 47254 20580 47292
rect 20636 47346 20692 47404
rect 20636 47294 20638 47346
rect 20690 47294 20692 47346
rect 20636 47236 20692 47294
rect 20636 47170 20692 47180
rect 20748 47068 20804 48076
rect 20748 47012 20916 47068
rect 20412 46386 20468 46396
rect 20636 46674 20692 46686
rect 20636 46622 20638 46674
rect 20690 46622 20692 46674
rect 20636 46116 20692 46622
rect 20860 46228 20916 47012
rect 20972 46786 21028 50764
rect 21084 50036 21140 50046
rect 21084 49942 21140 49980
rect 21196 49922 21252 49934
rect 21196 49870 21198 49922
rect 21250 49870 21252 49922
rect 21196 47572 21252 49870
rect 21308 49026 21364 52220
rect 21420 52274 21476 52332
rect 21420 52222 21422 52274
rect 21474 52222 21476 52274
rect 21420 52210 21476 52222
rect 21420 50372 21476 50382
rect 21420 50278 21476 50316
rect 21420 49812 21476 49822
rect 21532 49812 21588 54348
rect 22092 54290 22148 54302
rect 22092 54238 22094 54290
rect 22146 54238 22148 54290
rect 21756 53730 21812 53742
rect 21756 53678 21758 53730
rect 21810 53678 21812 53730
rect 21756 52948 21812 53678
rect 21420 49810 21588 49812
rect 21420 49758 21422 49810
rect 21474 49758 21588 49810
rect 21420 49756 21588 49758
rect 21644 52892 21756 52948
rect 21420 49746 21476 49756
rect 21308 48974 21310 49026
rect 21362 48974 21364 49026
rect 21308 48804 21364 48974
rect 21644 49028 21700 52892
rect 21756 52882 21812 52892
rect 21980 52948 22036 52958
rect 21868 52724 21924 52734
rect 21756 52722 21924 52724
rect 21756 52670 21870 52722
rect 21922 52670 21924 52722
rect 21756 52668 21924 52670
rect 21756 51268 21812 52668
rect 21868 52658 21924 52668
rect 21868 52164 21924 52174
rect 21868 52070 21924 52108
rect 21756 51202 21812 51212
rect 21868 50484 21924 50494
rect 21756 49812 21812 49822
rect 21756 49138 21812 49756
rect 21868 49810 21924 50428
rect 21868 49758 21870 49810
rect 21922 49758 21924 49810
rect 21868 49746 21924 49758
rect 21756 49086 21758 49138
rect 21810 49086 21812 49138
rect 21756 49074 21812 49086
rect 21868 49140 21924 49150
rect 21644 48934 21700 48972
rect 21868 49026 21924 49084
rect 21868 48974 21870 49026
rect 21922 48974 21924 49026
rect 21868 48962 21924 48974
rect 21308 48738 21364 48748
rect 21532 48916 21588 48926
rect 21532 48242 21588 48860
rect 21644 48468 21700 48478
rect 21644 48374 21700 48412
rect 21532 48190 21534 48242
rect 21586 48190 21588 48242
rect 21532 48178 21588 48190
rect 21196 47506 21252 47516
rect 21532 47460 21588 47470
rect 21532 47366 21588 47404
rect 20972 46734 20974 46786
rect 21026 46734 21028 46786
rect 20972 46722 21028 46734
rect 21196 47236 21252 47246
rect 21644 47236 21700 47246
rect 20860 46162 20916 46172
rect 20636 45892 20692 46060
rect 20188 45836 20468 45892
rect 20636 45836 21140 45892
rect 20076 45826 20132 45836
rect 19068 45666 19348 45668
rect 19068 45614 19070 45666
rect 19122 45614 19348 45666
rect 19068 45612 19348 45614
rect 19068 45602 19124 45612
rect 18956 45388 19236 45444
rect 18844 45332 18900 45342
rect 18844 45238 18900 45276
rect 19068 45220 19124 45230
rect 18956 45164 19068 45220
rect 18844 43764 18900 43774
rect 18788 43762 18900 43764
rect 18788 43710 18846 43762
rect 18898 43710 18900 43762
rect 18788 43708 18900 43710
rect 18732 43670 18788 43708
rect 18844 43698 18900 43708
rect 18732 43540 18788 43550
rect 18396 43426 18452 43438
rect 18396 43374 18398 43426
rect 18450 43374 18452 43426
rect 18396 43316 18452 43374
rect 18396 43250 18452 43260
rect 18732 43316 18788 43484
rect 18732 43250 18788 43260
rect 18844 42980 18900 42990
rect 18956 42980 19012 45164
rect 19068 45154 19124 45164
rect 19068 44324 19124 44334
rect 19068 43650 19124 44268
rect 19068 43598 19070 43650
rect 19122 43598 19124 43650
rect 19068 43586 19124 43598
rect 18844 42978 19012 42980
rect 18844 42926 18846 42978
rect 18898 42926 19012 42978
rect 18844 42924 19012 42926
rect 18844 42914 18900 42924
rect 18172 42754 18228 42812
rect 18172 42702 18174 42754
rect 18226 42702 18228 42754
rect 18172 42690 18228 42702
rect 18284 42756 18340 42766
rect 18284 42308 18340 42700
rect 18844 42756 18900 42766
rect 18284 42194 18340 42252
rect 18284 42142 18286 42194
rect 18338 42142 18340 42194
rect 18284 42130 18340 42142
rect 18732 42308 18788 42318
rect 18732 42082 18788 42252
rect 18844 42194 18900 42700
rect 18956 42754 19012 42766
rect 18956 42702 18958 42754
rect 19010 42702 19012 42754
rect 18956 42308 19012 42702
rect 18956 42242 19012 42252
rect 19068 42756 19124 42766
rect 18844 42142 18846 42194
rect 18898 42142 18900 42194
rect 18844 42130 18900 42142
rect 18732 42030 18734 42082
rect 18786 42030 18788 42082
rect 18732 42018 18788 42030
rect 19068 42084 19124 42700
rect 19180 42196 19236 45388
rect 19292 43876 19348 45612
rect 19516 45668 19572 45678
rect 19516 45574 19572 45612
rect 20300 45668 20356 45678
rect 20300 45574 20356 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19964 45218 20020 45230
rect 19964 45166 19966 45218
rect 20018 45166 20020 45218
rect 19852 45108 19908 45118
rect 19852 45014 19908 45052
rect 19964 44884 20020 45166
rect 19964 44818 20020 44828
rect 20188 45106 20244 45118
rect 20188 45054 20190 45106
rect 20242 45054 20244 45106
rect 19292 43810 19348 43820
rect 19516 44324 19572 44334
rect 19516 43538 19572 44268
rect 19628 44210 19684 44222
rect 19628 44158 19630 44210
rect 19682 44158 19684 44210
rect 19628 44100 19684 44158
rect 19628 44034 19684 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19516 43486 19518 43538
rect 19570 43486 19572 43538
rect 19516 43474 19572 43486
rect 19292 43428 19348 43438
rect 19292 43334 19348 43372
rect 19628 43428 19684 43438
rect 20188 43428 20244 45054
rect 20300 43428 20356 43438
rect 19684 43372 19796 43428
rect 20188 43426 20356 43428
rect 20188 43374 20302 43426
rect 20354 43374 20356 43426
rect 20188 43372 20356 43374
rect 19628 43362 19684 43372
rect 19628 42756 19684 42766
rect 19740 42756 19796 43372
rect 20300 43362 20356 43372
rect 19852 43316 19908 43326
rect 19852 43222 19908 43260
rect 19852 42756 19908 42766
rect 19740 42754 19908 42756
rect 19740 42702 19854 42754
rect 19906 42702 19908 42754
rect 19740 42700 19908 42702
rect 19628 42662 19684 42700
rect 19852 42690 19908 42700
rect 20300 42754 20356 42766
rect 20300 42702 20302 42754
rect 20354 42702 20356 42754
rect 20300 42644 20356 42702
rect 20300 42578 20356 42588
rect 19740 42532 19796 42570
rect 19740 42466 19796 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19180 42140 19796 42196
rect 19068 42028 19348 42084
rect 18396 41972 18452 41982
rect 18060 41916 18340 41972
rect 18060 41748 18116 41758
rect 18060 41746 18228 41748
rect 18060 41694 18062 41746
rect 18114 41694 18228 41746
rect 18060 41692 18228 41694
rect 18060 41682 18116 41692
rect 18060 40964 18116 40974
rect 17724 40516 17780 40526
rect 17948 40516 18004 40526
rect 17724 40422 17780 40460
rect 17836 40460 17948 40516
rect 17612 39442 17668 39452
rect 17836 39506 17892 40460
rect 17948 40450 18004 40460
rect 18060 40514 18116 40908
rect 18060 40462 18062 40514
rect 18114 40462 18116 40514
rect 18060 40450 18116 40462
rect 18060 40180 18116 40190
rect 18172 40180 18228 41692
rect 18284 41412 18340 41916
rect 18396 41858 18452 41916
rect 18396 41806 18398 41858
rect 18450 41806 18452 41858
rect 18396 41794 18452 41806
rect 19180 41860 19236 41870
rect 18844 41748 18900 41758
rect 18844 41746 19124 41748
rect 18844 41694 18846 41746
rect 18898 41694 19124 41746
rect 18844 41692 19124 41694
rect 18844 41682 18900 41692
rect 18284 41298 18340 41356
rect 18844 41412 18900 41422
rect 18844 41318 18900 41356
rect 18284 41246 18286 41298
rect 18338 41246 18340 41298
rect 18284 41234 18340 41246
rect 18620 41186 18676 41198
rect 18620 41134 18622 41186
rect 18674 41134 18676 41186
rect 18396 41076 18452 41086
rect 18284 40516 18340 40526
rect 18396 40516 18452 41020
rect 18620 40964 18676 41134
rect 18620 40898 18676 40908
rect 18284 40514 18452 40516
rect 18284 40462 18286 40514
rect 18338 40462 18452 40514
rect 18284 40460 18452 40462
rect 18732 40516 18788 40526
rect 18284 40450 18340 40460
rect 18732 40422 18788 40460
rect 18116 40124 18228 40180
rect 18396 40290 18452 40302
rect 18396 40238 18398 40290
rect 18450 40238 18452 40290
rect 18060 40114 18116 40124
rect 17836 39454 17838 39506
rect 17890 39454 17892 39506
rect 17836 39442 17892 39454
rect 18060 39618 18116 39630
rect 18060 39566 18062 39618
rect 18114 39566 18116 39618
rect 18060 39172 18116 39566
rect 18396 39620 18452 40238
rect 18956 40290 19012 40302
rect 18956 40238 18958 40290
rect 19010 40238 19012 40290
rect 18956 40180 19012 40238
rect 18956 40114 19012 40124
rect 19068 39620 19124 41692
rect 19180 41410 19236 41804
rect 19180 41358 19182 41410
rect 19234 41358 19236 41410
rect 19180 41346 19236 41358
rect 19180 40402 19236 40414
rect 19180 40350 19182 40402
rect 19234 40350 19236 40402
rect 19180 40068 19236 40350
rect 19180 40002 19236 40012
rect 19180 39620 19236 39630
rect 19068 39618 19236 39620
rect 19068 39566 19182 39618
rect 19234 39566 19236 39618
rect 19068 39564 19236 39566
rect 18396 39554 18452 39564
rect 19180 39554 19236 39564
rect 18956 39508 19012 39518
rect 18956 39414 19012 39452
rect 17388 39006 17390 39058
rect 17442 39006 17444 39058
rect 17388 38994 17444 39006
rect 17724 39116 18116 39172
rect 18732 39284 18788 39294
rect 17724 39058 17780 39116
rect 17724 39006 17726 39058
rect 17778 39006 17780 39058
rect 17276 38948 17332 38958
rect 17276 38668 17332 38892
rect 17724 38668 17780 39006
rect 17276 38612 17444 38668
rect 17164 37958 17220 37996
rect 17388 37938 17444 38612
rect 17388 37886 17390 37938
rect 17442 37886 17444 37938
rect 17388 36482 17444 37886
rect 17388 36430 17390 36482
rect 17442 36430 17444 36482
rect 17388 36418 17444 36430
rect 17500 38612 17780 38668
rect 18284 39060 18340 39070
rect 17500 37156 17556 38612
rect 18060 37716 18116 37726
rect 18060 37490 18116 37660
rect 18060 37438 18062 37490
rect 18114 37438 18116 37490
rect 18060 37426 18116 37438
rect 18172 37268 18228 37278
rect 18284 37268 18340 39004
rect 18508 39060 18564 39070
rect 18396 38836 18452 38846
rect 18396 37492 18452 38780
rect 18508 37716 18564 39004
rect 18508 37650 18564 37660
rect 18620 37492 18676 37502
rect 18396 37436 18564 37492
rect 18172 37266 18340 37268
rect 18172 37214 18174 37266
rect 18226 37214 18340 37266
rect 18172 37212 18340 37214
rect 18172 37202 18228 37212
rect 17388 36148 17444 36158
rect 17388 35138 17444 36092
rect 17388 35086 17390 35138
rect 17442 35086 17444 35138
rect 17388 35074 17444 35086
rect 17500 35586 17556 37100
rect 17724 37044 17780 37054
rect 18508 37044 18564 37436
rect 17612 36708 17668 36718
rect 17612 36614 17668 36652
rect 17724 35698 17780 36988
rect 17724 35646 17726 35698
rect 17778 35646 17780 35698
rect 17724 35634 17780 35646
rect 18172 36988 18564 37044
rect 17500 35534 17502 35586
rect 17554 35534 17556 35586
rect 17052 33516 17220 33572
rect 16604 33348 16660 33358
rect 16604 33254 16660 33292
rect 17052 33346 17108 33358
rect 17052 33294 17054 33346
rect 17106 33294 17108 33346
rect 17052 33236 17108 33294
rect 16492 33122 16548 33134
rect 16492 33070 16494 33122
rect 16546 33070 16548 33122
rect 16492 32676 16548 33070
rect 16492 32610 16548 32620
rect 16604 33012 16660 33022
rect 16380 31266 16436 31276
rect 15820 31220 15876 31230
rect 15820 30994 15876 31164
rect 15820 30942 15822 30994
rect 15874 30942 15876 30994
rect 15708 30884 15764 30894
rect 15596 30882 15764 30884
rect 15596 30830 15710 30882
rect 15762 30830 15764 30882
rect 15596 30828 15764 30830
rect 15708 30818 15764 30828
rect 14812 30156 15316 30212
rect 14924 29988 14980 29998
rect 14700 29986 14980 29988
rect 14700 29934 14926 29986
rect 14978 29934 14980 29986
rect 14700 29932 14980 29934
rect 14924 29922 14980 29932
rect 15260 29988 15316 30156
rect 15820 30210 15876 30942
rect 16604 30434 16660 32956
rect 17052 32564 17108 33180
rect 17052 32498 17108 32508
rect 17164 31892 17220 33516
rect 17276 33236 17332 33246
rect 17500 33236 17556 35534
rect 18060 35588 18116 35598
rect 18060 35494 18116 35532
rect 17836 35476 17892 35486
rect 17724 34356 17780 34366
rect 17724 34262 17780 34300
rect 17836 33458 17892 35420
rect 18060 35364 18116 35374
rect 17836 33406 17838 33458
rect 17890 33406 17892 33458
rect 17836 33394 17892 33406
rect 17948 34692 18004 34702
rect 17276 33234 17556 33236
rect 17276 33182 17278 33234
rect 17330 33182 17556 33234
rect 17276 33180 17556 33182
rect 17276 33170 17332 33180
rect 17836 32900 17892 32910
rect 17836 32562 17892 32844
rect 17836 32510 17838 32562
rect 17890 32510 17892 32562
rect 17836 32498 17892 32510
rect 17948 32788 18004 34636
rect 18060 33458 18116 35308
rect 18172 34132 18228 36988
rect 18396 36820 18452 36830
rect 18396 35026 18452 36764
rect 18620 36708 18676 37436
rect 18508 36652 18676 36708
rect 18508 35924 18564 36652
rect 18732 36594 18788 39228
rect 19068 39284 19124 39294
rect 18844 37604 18900 37614
rect 18844 37044 18900 37548
rect 18956 37492 19012 37502
rect 18956 37378 19012 37436
rect 18956 37326 18958 37378
rect 19010 37326 19012 37378
rect 18956 37314 19012 37326
rect 18844 36978 18900 36988
rect 18956 36820 19012 36830
rect 18732 36542 18734 36594
rect 18786 36542 18788 36594
rect 18620 36484 18676 36494
rect 18620 36390 18676 36428
rect 18508 35868 18676 35924
rect 18508 35700 18564 35710
rect 18508 35606 18564 35644
rect 18620 35252 18676 35868
rect 18396 34974 18398 35026
rect 18450 34974 18452 35026
rect 18396 34962 18452 34974
rect 18508 35196 18676 35252
rect 18284 34132 18340 34142
rect 18172 34130 18340 34132
rect 18172 34078 18286 34130
rect 18338 34078 18340 34130
rect 18172 34076 18340 34078
rect 18284 34066 18340 34076
rect 18060 33406 18062 33458
rect 18114 33406 18116 33458
rect 18060 33394 18116 33406
rect 18508 33346 18564 35196
rect 18620 34804 18676 34814
rect 18620 34130 18676 34748
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18620 34066 18676 34078
rect 18508 33294 18510 33346
rect 18562 33294 18564 33346
rect 18508 33124 18564 33294
rect 18620 33458 18676 33470
rect 18620 33406 18622 33458
rect 18674 33406 18676 33458
rect 18620 33236 18676 33406
rect 18620 33170 18676 33180
rect 18508 33058 18564 33068
rect 17948 32450 18004 32732
rect 18732 32564 18788 36542
rect 18844 36596 18900 36606
rect 18844 36372 18900 36540
rect 18956 36594 19012 36764
rect 18956 36542 18958 36594
rect 19010 36542 19012 36594
rect 18956 36530 19012 36542
rect 18844 36316 19012 36372
rect 18844 34356 18900 34366
rect 18844 34130 18900 34300
rect 18844 34078 18846 34130
rect 18898 34078 18900 34130
rect 18844 34066 18900 34078
rect 18844 33572 18900 33582
rect 18844 33012 18900 33516
rect 18844 32946 18900 32956
rect 18956 32788 19012 36316
rect 19068 34356 19124 39228
rect 19292 38668 19348 42028
rect 19516 41074 19572 41086
rect 19516 41022 19518 41074
rect 19570 41022 19572 41074
rect 19516 40964 19572 41022
rect 19740 41076 19796 42140
rect 19852 42084 19908 42094
rect 20412 42084 20468 45836
rect 20748 45668 20804 45678
rect 20524 45666 20804 45668
rect 20524 45614 20750 45666
rect 20802 45614 20804 45666
rect 20524 45612 20804 45614
rect 20524 44548 20580 45612
rect 20748 45602 20804 45612
rect 20524 44482 20580 44492
rect 20748 44324 20804 44334
rect 20748 44322 20916 44324
rect 20748 44270 20750 44322
rect 20802 44270 20916 44322
rect 20748 44268 20916 44270
rect 20748 44258 20804 44268
rect 20524 44098 20580 44110
rect 20524 44046 20526 44098
rect 20578 44046 20580 44098
rect 20524 43538 20580 44046
rect 20860 43652 20916 44268
rect 20972 43652 21028 43662
rect 20860 43596 20972 43652
rect 20972 43586 21028 43596
rect 20524 43486 20526 43538
rect 20578 43486 20580 43538
rect 20524 43474 20580 43486
rect 20524 42642 20580 42654
rect 20524 42590 20526 42642
rect 20578 42590 20580 42642
rect 20524 42308 20580 42590
rect 20636 42532 20692 42542
rect 20636 42438 20692 42476
rect 20860 42532 20916 42542
rect 20860 42438 20916 42476
rect 20524 42242 20580 42252
rect 20972 42308 21028 42318
rect 20412 42028 20692 42084
rect 19852 41858 19908 42028
rect 19852 41806 19854 41858
rect 19906 41806 19908 41858
rect 19852 41794 19908 41806
rect 19964 41858 20020 41870
rect 19964 41806 19966 41858
rect 20018 41806 20020 41858
rect 19964 41412 20020 41806
rect 19964 41346 20020 41356
rect 20412 41858 20468 41870
rect 20412 41806 20414 41858
rect 20466 41806 20468 41858
rect 20412 41748 20468 41806
rect 19740 40982 19796 41020
rect 19516 40898 19572 40908
rect 19628 40962 19684 40974
rect 19628 40910 19630 40962
rect 19682 40910 19684 40962
rect 19628 40628 19684 40910
rect 20300 40964 20356 40974
rect 20300 40870 20356 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40572 20132 40628
rect 20076 40570 20132 40572
rect 20076 40518 20078 40570
rect 20130 40518 20132 40570
rect 20076 40506 20132 40518
rect 19852 40404 19908 40414
rect 19628 40348 19852 40404
rect 19516 40068 19572 40078
rect 19404 39956 19460 39966
rect 19404 39730 19460 39900
rect 19404 39678 19406 39730
rect 19458 39678 19460 39730
rect 19404 39666 19460 39678
rect 19516 39506 19572 40012
rect 19516 39454 19518 39506
rect 19570 39454 19572 39506
rect 19516 38836 19572 39454
rect 19628 39060 19684 40348
rect 19852 40310 19908 40348
rect 20300 40402 20356 40414
rect 20300 40350 20302 40402
rect 20354 40350 20356 40402
rect 20188 40290 20244 40302
rect 20188 40238 20190 40290
rect 20242 40238 20244 40290
rect 19964 40180 20020 40190
rect 19964 39732 20020 40124
rect 19964 39638 20020 39676
rect 20188 39618 20244 40238
rect 20300 40180 20356 40350
rect 20300 40114 20356 40124
rect 20188 39566 20190 39618
rect 20242 39566 20244 39618
rect 20188 39554 20244 39566
rect 20412 39396 20468 41692
rect 20636 40964 20692 42028
rect 20972 41858 21028 42252
rect 20972 41806 20974 41858
rect 21026 41806 21028 41858
rect 20972 41636 21028 41806
rect 20972 41570 21028 41580
rect 20748 40964 20804 40974
rect 20524 40962 20804 40964
rect 20524 40910 20750 40962
rect 20802 40910 20804 40962
rect 20524 40908 20804 40910
rect 20524 40404 20580 40908
rect 20748 40898 20804 40908
rect 20748 40740 20804 40750
rect 20524 40338 20580 40348
rect 20636 40402 20692 40414
rect 20636 40350 20638 40402
rect 20690 40350 20692 40402
rect 20636 40292 20692 40350
rect 20636 40226 20692 40236
rect 20524 39620 20580 39630
rect 20524 39526 20580 39564
rect 20412 39330 20468 39340
rect 20748 39506 20804 40684
rect 20748 39454 20750 39506
rect 20802 39454 20804 39506
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19628 39004 20020 39060
rect 19628 38836 19684 38846
rect 19516 38780 19628 38836
rect 19628 38770 19684 38780
rect 19964 38834 20020 39004
rect 20748 38948 20804 39454
rect 20860 39396 20916 39406
rect 20860 39394 21028 39396
rect 20860 39342 20862 39394
rect 20914 39342 21028 39394
rect 20860 39340 21028 39342
rect 20860 39330 20916 39340
rect 20860 38948 20916 38958
rect 20748 38946 20916 38948
rect 20748 38894 20862 38946
rect 20914 38894 20916 38946
rect 20748 38892 20916 38894
rect 20860 38882 20916 38892
rect 19964 38782 19966 38834
rect 20018 38782 20020 38834
rect 19964 38770 20020 38782
rect 20412 38834 20468 38846
rect 20412 38782 20414 38834
rect 20466 38782 20468 38834
rect 20412 38668 20468 38782
rect 19292 38612 19684 38668
rect 19292 38164 19348 38174
rect 19292 38050 19348 38108
rect 19292 37998 19294 38050
rect 19346 37998 19348 38050
rect 19292 37986 19348 37998
rect 19516 38050 19572 38062
rect 19516 37998 19518 38050
rect 19570 37998 19572 38050
rect 19516 37492 19572 37998
rect 19628 37938 19684 38612
rect 20300 38612 20468 38668
rect 19628 37886 19630 37938
rect 19682 37886 19684 37938
rect 19628 37492 19684 37886
rect 19740 38164 19796 38174
rect 19740 37940 19796 38108
rect 19740 37874 19796 37884
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37436 20244 37492
rect 19516 37426 19572 37436
rect 19292 37268 19348 37278
rect 19292 36482 19348 37212
rect 19516 37268 19572 37278
rect 19292 36430 19294 36482
rect 19346 36430 19348 36482
rect 19292 36418 19348 36430
rect 19404 36484 19460 36494
rect 19404 35698 19460 36428
rect 19404 35646 19406 35698
rect 19458 35646 19460 35698
rect 19292 35476 19348 35486
rect 19180 35252 19236 35262
rect 19180 34804 19236 35196
rect 19292 34914 19348 35420
rect 19404 35138 19460 35646
rect 19404 35086 19406 35138
rect 19458 35086 19460 35138
rect 19404 35074 19460 35086
rect 19516 36370 19572 37212
rect 19852 37266 19908 37278
rect 19852 37214 19854 37266
rect 19906 37214 19908 37266
rect 19852 37156 19908 37214
rect 19852 37090 19908 37100
rect 19516 36318 19518 36370
rect 19570 36318 19572 36370
rect 19292 34862 19294 34914
rect 19346 34862 19348 34914
rect 19292 34850 19348 34862
rect 19180 34710 19236 34748
rect 19180 34356 19236 34366
rect 19068 34354 19236 34356
rect 19068 34302 19182 34354
rect 19234 34302 19236 34354
rect 19068 34300 19236 34302
rect 19180 34290 19236 34300
rect 19516 34132 19572 36318
rect 18956 32722 19012 32732
rect 19068 34076 19572 34132
rect 19628 37044 19684 37054
rect 19068 32674 19124 34076
rect 19628 34020 19684 36988
rect 20076 36594 20132 36606
rect 20076 36542 20078 36594
rect 20130 36542 20132 36594
rect 20076 36372 20132 36542
rect 20188 36482 20244 37436
rect 20300 37044 20356 38612
rect 20412 38546 20468 38556
rect 20972 38276 21028 39340
rect 21084 39060 21140 45836
rect 21196 40964 21252 47180
rect 21532 47180 21644 47236
rect 21308 47124 21364 47134
rect 21308 46788 21364 47068
rect 21308 46694 21364 46732
rect 21420 46786 21476 46798
rect 21420 46734 21422 46786
rect 21474 46734 21476 46786
rect 21420 46564 21476 46734
rect 21308 44324 21364 44334
rect 21308 44230 21364 44268
rect 21308 42980 21364 42990
rect 21308 41748 21364 42924
rect 21420 42196 21476 46508
rect 21420 42130 21476 42140
rect 21420 41858 21476 41870
rect 21420 41806 21422 41858
rect 21474 41806 21476 41858
rect 21420 41748 21476 41806
rect 21308 41746 21476 41748
rect 21308 41694 21310 41746
rect 21362 41694 21476 41746
rect 21308 41692 21476 41694
rect 21308 41682 21364 41692
rect 21532 41636 21588 47180
rect 21644 47170 21700 47180
rect 21644 46676 21700 46686
rect 21868 46676 21924 46686
rect 21644 46674 21924 46676
rect 21644 46622 21646 46674
rect 21698 46622 21870 46674
rect 21922 46622 21924 46674
rect 21644 46620 21924 46622
rect 21644 46610 21700 46620
rect 21868 46610 21924 46620
rect 21980 46228 22036 52892
rect 22092 52946 22148 54238
rect 22652 54290 22708 54302
rect 22652 54238 22654 54290
rect 22706 54238 22708 54290
rect 22652 54180 22708 54238
rect 22652 54114 22708 54124
rect 22764 54290 22820 54796
rect 22764 54238 22766 54290
rect 22818 54238 22820 54290
rect 22764 53956 22820 54238
rect 22316 53900 22820 53956
rect 22876 54180 22932 55020
rect 23324 54516 23380 55020
rect 23324 54422 23380 54460
rect 23660 54628 23716 54638
rect 23772 54628 23828 55246
rect 24892 55186 24948 55198
rect 24892 55134 24894 55186
rect 24946 55134 24948 55186
rect 24892 54852 24948 55134
rect 24892 54786 24948 54796
rect 23716 54572 23828 54628
rect 23660 54514 23716 54572
rect 23660 54462 23662 54514
rect 23714 54462 23716 54514
rect 22316 53730 22372 53900
rect 22540 53732 22596 53742
rect 22316 53678 22318 53730
rect 22370 53678 22372 53730
rect 22316 53508 22372 53678
rect 22316 53442 22372 53452
rect 22428 53676 22540 53732
rect 22092 52894 22094 52946
rect 22146 52894 22148 52946
rect 22092 52882 22148 52894
rect 22316 52834 22372 52846
rect 22316 52782 22318 52834
rect 22370 52782 22372 52834
rect 22092 52276 22148 52286
rect 22092 52162 22148 52220
rect 22092 52110 22094 52162
rect 22146 52110 22148 52162
rect 22092 52098 22148 52110
rect 22316 52052 22372 52782
rect 22316 51986 22372 51996
rect 22428 51380 22484 53676
rect 22540 53638 22596 53676
rect 22876 53730 22932 54124
rect 22876 53678 22878 53730
rect 22930 53678 22932 53730
rect 22764 53172 22820 53182
rect 22764 53078 22820 53116
rect 22540 52948 22596 52958
rect 22540 52854 22596 52892
rect 22652 52834 22708 52846
rect 22652 52782 22654 52834
rect 22706 52782 22708 52834
rect 22652 52164 22708 52782
rect 22764 52164 22820 52174
rect 22652 52162 22820 52164
rect 22652 52110 22766 52162
rect 22818 52110 22820 52162
rect 22652 52108 22820 52110
rect 22764 52098 22820 52108
rect 22204 51324 22484 51380
rect 22540 51378 22596 51390
rect 22540 51326 22542 51378
rect 22594 51326 22596 51378
rect 22092 50596 22148 50634
rect 22092 50530 22148 50540
rect 22204 50428 22260 51324
rect 22540 51156 22596 51326
rect 22428 51100 22540 51156
rect 22316 50596 22372 50606
rect 22316 50502 22372 50540
rect 22092 50372 22260 50428
rect 22428 50428 22484 51100
rect 22540 51090 22596 51100
rect 22652 51380 22708 51390
rect 22540 50708 22596 50718
rect 22652 50708 22708 51324
rect 22876 50820 22932 53678
rect 23436 54290 23492 54302
rect 23436 54238 23438 54290
rect 23490 54238 23492 54290
rect 23436 54068 23492 54238
rect 23660 54068 23716 54462
rect 25116 54516 25172 56030
rect 25788 55972 25844 56252
rect 25788 55970 25956 55972
rect 25788 55918 25790 55970
rect 25842 55918 25956 55970
rect 25788 55916 25956 55918
rect 25788 55906 25844 55916
rect 25116 54450 25172 54460
rect 25228 55858 25284 55870
rect 25228 55806 25230 55858
rect 25282 55806 25284 55858
rect 23772 54292 23828 54302
rect 23772 54290 24836 54292
rect 23772 54238 23774 54290
rect 23826 54238 24836 54290
rect 23772 54236 24836 54238
rect 23772 54226 23828 54236
rect 23436 54012 23604 54068
rect 23660 54012 24052 54068
rect 23436 53732 23492 54012
rect 23548 53956 23604 54012
rect 23548 53900 23828 53956
rect 23772 53842 23828 53900
rect 23772 53790 23774 53842
rect 23826 53790 23828 53842
rect 23772 53778 23828 53790
rect 23884 53844 23940 53854
rect 23884 53750 23940 53788
rect 23436 53666 23492 53676
rect 23996 53618 24052 54012
rect 24780 53730 24836 54236
rect 25228 53844 25284 55806
rect 25676 55188 25732 55198
rect 25228 53778 25284 53788
rect 25340 55186 25732 55188
rect 25340 55134 25678 55186
rect 25730 55134 25732 55186
rect 25340 55132 25732 55134
rect 25116 53732 25172 53742
rect 24780 53678 24782 53730
rect 24834 53678 24836 53730
rect 24780 53666 24836 53678
rect 25004 53730 25172 53732
rect 25004 53678 25118 53730
rect 25170 53678 25172 53730
rect 25004 53676 25172 53678
rect 23996 53566 23998 53618
rect 24050 53566 24052 53618
rect 23996 53554 24052 53566
rect 23100 53506 23156 53518
rect 23100 53454 23102 53506
rect 23154 53454 23156 53506
rect 23100 53172 23156 53454
rect 22988 52388 23044 52398
rect 22988 52294 23044 52332
rect 23100 52276 23156 53116
rect 23324 53508 23380 53518
rect 23324 53170 23380 53452
rect 23324 53118 23326 53170
rect 23378 53118 23380 53170
rect 23212 52948 23268 52958
rect 23212 52388 23268 52892
rect 23212 52322 23268 52332
rect 23100 52210 23156 52220
rect 23324 52164 23380 53118
rect 23436 53284 23492 53294
rect 23436 52386 23492 53228
rect 24556 52836 24612 52846
rect 23436 52334 23438 52386
rect 23490 52334 23492 52386
rect 23436 52322 23492 52334
rect 24444 52834 24612 52836
rect 24444 52782 24558 52834
rect 24610 52782 24612 52834
rect 24444 52780 24612 52782
rect 23660 52164 23716 52174
rect 23324 52162 23716 52164
rect 23324 52110 23662 52162
rect 23714 52110 23716 52162
rect 23324 52108 23716 52110
rect 23660 52098 23716 52108
rect 23996 52164 24052 52174
rect 23996 52070 24052 52108
rect 23772 52052 23828 52062
rect 22988 51604 23044 51614
rect 23772 51604 23828 51996
rect 23884 51940 23940 51950
rect 23884 51846 23940 51884
rect 24108 51940 24164 51950
rect 24444 51940 24500 52780
rect 24556 52770 24612 52780
rect 25004 52276 25060 53676
rect 25116 53666 25172 53676
rect 25116 53506 25172 53518
rect 25116 53454 25118 53506
rect 25170 53454 25172 53506
rect 25116 53172 25172 53454
rect 25340 53284 25396 55132
rect 25676 55122 25732 55132
rect 25788 55074 25844 55086
rect 25788 55022 25790 55074
rect 25842 55022 25844 55074
rect 25788 54628 25844 55022
rect 25900 54852 25956 55916
rect 26908 55970 26964 55982
rect 26908 55918 26910 55970
rect 26962 55918 26964 55970
rect 26908 55468 26964 55918
rect 29596 55970 29652 59200
rect 34300 56308 34356 56318
rect 33740 56306 34356 56308
rect 33740 56254 34302 56306
rect 34354 56254 34356 56306
rect 33740 56252 34356 56254
rect 33740 56194 33796 56252
rect 34300 56242 34356 56252
rect 47740 56308 47796 59200
rect 47740 56242 47796 56252
rect 33740 56142 33742 56194
rect 33794 56142 33796 56194
rect 31164 56084 31220 56094
rect 31164 55990 31220 56028
rect 32284 56084 32340 56094
rect 32284 55990 32340 56028
rect 33292 56082 33348 56094
rect 33292 56030 33294 56082
rect 33346 56030 33348 56082
rect 29596 55918 29598 55970
rect 29650 55918 29652 55970
rect 29596 55906 29652 55918
rect 26684 55412 26964 55468
rect 31612 55748 31668 55758
rect 29372 55412 29428 55422
rect 26460 55186 26516 55198
rect 26460 55134 26462 55186
rect 26514 55134 26516 55186
rect 26012 55076 26068 55086
rect 26012 55074 26404 55076
rect 26012 55022 26014 55074
rect 26066 55022 26404 55074
rect 26012 55020 26404 55022
rect 26012 55010 26068 55020
rect 25900 54796 26068 54852
rect 25340 53218 25396 53228
rect 25452 54572 25844 54628
rect 25452 53618 25508 54572
rect 25900 54516 25956 54554
rect 25900 54450 25956 54460
rect 25676 54404 25732 54414
rect 25676 54310 25732 54348
rect 25564 54292 25620 54302
rect 25564 53956 25620 54236
rect 25564 53890 25620 53900
rect 25788 53844 25844 53854
rect 25788 53730 25844 53788
rect 25788 53678 25790 53730
rect 25842 53678 25844 53730
rect 25788 53666 25844 53678
rect 25452 53566 25454 53618
rect 25506 53566 25508 53618
rect 25116 53106 25172 53116
rect 25340 52276 25396 52314
rect 25004 52220 25172 52276
rect 24108 51938 24500 51940
rect 24108 51886 24110 51938
rect 24162 51886 24500 51938
rect 24108 51884 24500 51886
rect 24556 52162 24612 52174
rect 24556 52110 24558 52162
rect 24610 52110 24612 52162
rect 24108 51874 24164 51884
rect 23884 51604 23940 51614
rect 23772 51548 23884 51604
rect 22988 51510 23044 51548
rect 23884 51510 23940 51548
rect 23212 51490 23268 51502
rect 23212 51438 23214 51490
rect 23266 51438 23268 51490
rect 23212 51044 23268 51438
rect 23660 51492 23716 51502
rect 23660 51398 23716 51436
rect 24108 51380 24164 51390
rect 24108 51286 24164 51324
rect 23996 51266 24052 51278
rect 23996 51214 23998 51266
rect 24050 51214 24052 51266
rect 23212 50978 23268 50988
rect 23884 51156 23940 51166
rect 22876 50764 23268 50820
rect 22540 50706 22708 50708
rect 22540 50654 22542 50706
rect 22594 50654 22708 50706
rect 22540 50652 22708 50654
rect 22540 50642 22596 50652
rect 23212 50596 23268 50764
rect 23884 50706 23940 51100
rect 23996 50820 24052 51214
rect 24220 51156 24276 51884
rect 24556 51602 24612 52110
rect 25004 52050 25060 52062
rect 25004 51998 25006 52050
rect 25058 51998 25060 52050
rect 25004 51940 25060 51998
rect 24556 51550 24558 51602
rect 24610 51550 24612 51602
rect 24332 51156 24388 51166
rect 24220 51154 24388 51156
rect 24220 51102 24334 51154
rect 24386 51102 24388 51154
rect 24220 51100 24388 51102
rect 24332 51090 24388 51100
rect 23996 50764 24388 50820
rect 23884 50654 23886 50706
rect 23938 50654 23940 50706
rect 23884 50642 23940 50654
rect 23212 50530 23268 50540
rect 23996 50596 24052 50606
rect 22652 50484 22708 50494
rect 22988 50484 23044 50494
rect 22428 50372 22708 50428
rect 22764 50482 23044 50484
rect 22764 50430 22990 50482
rect 23042 50430 23044 50482
rect 22764 50428 23044 50430
rect 22092 46452 22148 50372
rect 22764 50036 22820 50428
rect 22988 50418 23044 50428
rect 23100 50484 23156 50522
rect 23772 50482 23828 50494
rect 23772 50430 23774 50482
rect 23826 50430 23828 50482
rect 23772 50428 23828 50430
rect 23100 50418 23156 50428
rect 23324 50372 23380 50382
rect 22428 49980 22820 50036
rect 23212 50370 23380 50372
rect 23212 50318 23326 50370
rect 23378 50318 23380 50370
rect 23212 50316 23380 50318
rect 22428 49812 22484 49980
rect 22652 49812 22708 49822
rect 22428 49746 22484 49756
rect 22540 49756 22652 49812
rect 22428 49588 22484 49598
rect 22204 48802 22260 48814
rect 22204 48750 22206 48802
rect 22258 48750 22260 48802
rect 22204 47236 22260 48750
rect 22204 47170 22260 47180
rect 22316 48020 22372 48030
rect 22316 47570 22372 47964
rect 22316 47518 22318 47570
rect 22370 47518 22372 47570
rect 22092 46386 22148 46396
rect 21980 46172 22260 46228
rect 21868 45892 21924 45902
rect 21868 44548 21924 45836
rect 22204 45332 22260 46172
rect 22092 44996 22148 45006
rect 22092 44902 22148 44940
rect 21868 44482 21924 44492
rect 21756 44324 21812 44334
rect 21756 44230 21812 44268
rect 22092 44210 22148 44222
rect 22092 44158 22094 44210
rect 22146 44158 22148 44210
rect 22092 44100 22148 44158
rect 22092 44034 22148 44044
rect 21756 43876 21812 43886
rect 21756 43314 21812 43820
rect 22204 43538 22260 45276
rect 22204 43486 22206 43538
rect 22258 43486 22260 43538
rect 22204 43474 22260 43486
rect 21756 43262 21758 43314
rect 21810 43262 21812 43314
rect 21756 43250 21812 43262
rect 21644 42868 21700 42878
rect 21644 42774 21700 42812
rect 21756 42756 21812 42766
rect 21980 42756 22036 42766
rect 21756 42662 21812 42700
rect 21868 42754 22036 42756
rect 21868 42702 21982 42754
rect 22034 42702 22036 42754
rect 21868 42700 22036 42702
rect 21644 42196 21700 42206
rect 21644 42102 21700 42140
rect 21196 40402 21252 40908
rect 21196 40350 21198 40402
rect 21250 40350 21252 40402
rect 21196 40338 21252 40350
rect 21420 41580 21588 41636
rect 21420 39732 21476 41580
rect 21532 41412 21588 41422
rect 21868 41412 21924 42700
rect 21980 42690 22036 42700
rect 21588 41356 21924 41412
rect 21980 41970 22036 41982
rect 21980 41918 21982 41970
rect 22034 41918 22036 41970
rect 21532 41298 21588 41356
rect 21532 41246 21534 41298
rect 21586 41246 21588 41298
rect 21532 41076 21588 41246
rect 21532 41010 21588 41020
rect 21980 41300 22036 41918
rect 22316 41412 22372 47518
rect 22428 46676 22484 49532
rect 22540 48914 22596 49756
rect 22652 49746 22708 49756
rect 23212 49810 23268 50316
rect 23324 50306 23380 50316
rect 23660 50372 23828 50428
rect 23660 50148 23716 50372
rect 23996 50370 24052 50540
rect 23996 50318 23998 50370
rect 24050 50318 24052 50370
rect 23996 50306 24052 50318
rect 23660 50092 24052 50148
rect 23772 49812 23828 50092
rect 23212 49758 23214 49810
rect 23266 49758 23268 49810
rect 23212 49746 23268 49758
rect 23548 49756 23828 49812
rect 23548 49698 23604 49756
rect 23548 49646 23550 49698
rect 23602 49646 23604 49698
rect 23548 49634 23604 49646
rect 22988 49588 23044 49598
rect 22988 49494 23044 49532
rect 23772 49588 23828 49598
rect 23212 49252 23268 49262
rect 23268 49196 23380 49252
rect 23212 49186 23268 49196
rect 22540 48862 22542 48914
rect 22594 48862 22596 48914
rect 22540 48850 22596 48862
rect 22876 49028 22932 49038
rect 22876 48914 22932 48972
rect 22876 48862 22878 48914
rect 22930 48862 22932 48914
rect 22876 48850 22932 48862
rect 23212 48804 23268 48814
rect 23212 48710 23268 48748
rect 22540 48692 22596 48702
rect 22540 47460 22596 48636
rect 23324 48466 23380 49196
rect 23772 49026 23828 49532
rect 23884 49586 23940 49598
rect 23884 49534 23886 49586
rect 23938 49534 23940 49586
rect 23884 49252 23940 49534
rect 23884 49186 23940 49196
rect 23996 49028 24052 50092
rect 24108 49922 24164 49934
rect 24108 49870 24110 49922
rect 24162 49870 24164 49922
rect 24108 49812 24164 49870
rect 24108 49746 24164 49756
rect 24220 49700 24276 49710
rect 24220 49606 24276 49644
rect 23772 48974 23774 49026
rect 23826 48974 23828 49026
rect 23772 48962 23828 48974
rect 23884 48972 24052 49028
rect 23324 48414 23326 48466
rect 23378 48414 23380 48466
rect 23324 48402 23380 48414
rect 23548 48914 23604 48926
rect 23548 48862 23550 48914
rect 23602 48862 23604 48914
rect 22652 48354 22708 48366
rect 22652 48302 22654 48354
rect 22706 48302 22708 48354
rect 22652 48244 22708 48302
rect 22652 48178 22708 48188
rect 23548 48244 23604 48862
rect 23548 48178 23604 48188
rect 23212 48018 23268 48030
rect 23212 47966 23214 48018
rect 23266 47966 23268 48018
rect 23212 47908 23268 47966
rect 23548 48020 23604 48030
rect 23548 47926 23604 47964
rect 22988 47852 23268 47908
rect 22764 47572 22820 47582
rect 22596 47404 22708 47460
rect 22540 47366 22596 47404
rect 22540 46676 22596 46686
rect 22428 46674 22596 46676
rect 22428 46622 22542 46674
rect 22594 46622 22596 46674
rect 22428 46620 22596 46622
rect 22540 46452 22596 46620
rect 22540 46386 22596 46396
rect 22652 46562 22708 47404
rect 22764 47234 22820 47516
rect 22988 47570 23044 47852
rect 22988 47518 22990 47570
rect 23042 47518 23044 47570
rect 22764 47182 22766 47234
rect 22818 47182 22820 47234
rect 22764 47170 22820 47182
rect 22876 47236 22932 47246
rect 22876 47142 22932 47180
rect 22988 46788 23044 47518
rect 23548 47348 23604 47358
rect 23548 47346 23716 47348
rect 23548 47294 23550 47346
rect 23602 47294 23716 47346
rect 23548 47292 23716 47294
rect 23548 47282 23604 47292
rect 23324 47236 23380 47246
rect 23324 47142 23380 47180
rect 23436 47234 23492 47246
rect 23436 47182 23438 47234
rect 23490 47182 23492 47234
rect 23436 47012 23492 47182
rect 23548 47124 23604 47134
rect 23660 47124 23716 47292
rect 23884 47236 23940 48972
rect 24332 48804 24388 50764
rect 24332 48738 24388 48748
rect 24556 48692 24612 51550
rect 24892 51604 24948 51614
rect 24892 51268 24948 51548
rect 25004 51492 25060 51884
rect 25116 51604 25172 52220
rect 25340 52210 25396 52220
rect 25340 52052 25396 52062
rect 25340 51958 25396 51996
rect 25116 51548 25284 51604
rect 25004 51426 25060 51436
rect 25116 51378 25172 51390
rect 25116 51326 25118 51378
rect 25170 51326 25172 51378
rect 25004 51268 25060 51278
rect 24892 51212 25004 51268
rect 24780 51154 24836 51166
rect 24780 51102 24782 51154
rect 24834 51102 24836 51154
rect 24780 50428 24836 51102
rect 25004 50482 25060 51212
rect 25004 50430 25006 50482
rect 25058 50430 25060 50482
rect 24780 50372 24948 50428
rect 25004 50418 25060 50430
rect 24668 49698 24724 49710
rect 24668 49646 24670 49698
rect 24722 49646 24724 49698
rect 24668 49476 24724 49646
rect 24668 49410 24724 49420
rect 24556 48626 24612 48636
rect 24108 48130 24164 48142
rect 24780 48132 24836 48142
rect 24108 48078 24110 48130
rect 24162 48078 24164 48130
rect 24108 47796 24164 48078
rect 24668 48130 24836 48132
rect 24668 48078 24782 48130
rect 24834 48078 24836 48130
rect 24668 48076 24836 48078
rect 24668 48020 24724 48076
rect 24780 48066 24836 48076
rect 24108 47740 24500 47796
rect 24332 47572 24388 47582
rect 23996 47570 24388 47572
rect 23996 47518 24334 47570
rect 24386 47518 24388 47570
rect 23996 47516 24388 47518
rect 23996 47458 24052 47516
rect 24332 47506 24388 47516
rect 23996 47406 23998 47458
rect 24050 47406 24052 47458
rect 23996 47394 24052 47406
rect 24444 47458 24500 47740
rect 24444 47406 24446 47458
rect 24498 47406 24500 47458
rect 24220 47346 24276 47358
rect 24220 47294 24222 47346
rect 24274 47294 24276 47346
rect 24108 47236 24164 47246
rect 23884 47180 24052 47236
rect 23604 47068 23716 47124
rect 23548 47058 23604 47068
rect 23436 46946 23492 46956
rect 23324 46900 23380 46910
rect 22988 46722 23044 46732
rect 23100 46786 23156 46798
rect 23100 46734 23102 46786
rect 23154 46734 23156 46786
rect 22652 46510 22654 46562
rect 22706 46510 22708 46562
rect 22428 46340 22484 46350
rect 22428 44434 22484 46284
rect 22652 45388 22708 46510
rect 23100 46116 23156 46734
rect 23100 46050 23156 46060
rect 23100 45890 23156 45902
rect 23100 45838 23102 45890
rect 23154 45838 23156 45890
rect 22652 45332 22932 45388
rect 22428 44382 22430 44434
rect 22482 44382 22484 44434
rect 22428 44324 22484 44382
rect 22428 44258 22484 44268
rect 22540 45108 22596 45118
rect 22540 42866 22596 45052
rect 22764 45106 22820 45118
rect 22764 45054 22766 45106
rect 22818 45054 22820 45106
rect 22652 44996 22708 45006
rect 22652 44902 22708 44940
rect 22764 44660 22820 45054
rect 22764 44594 22820 44604
rect 22652 44212 22708 44222
rect 22708 44156 22820 44212
rect 22652 44146 22708 44156
rect 22540 42814 22542 42866
rect 22594 42814 22596 42866
rect 22540 42802 22596 42814
rect 22652 41972 22708 41982
rect 22652 41878 22708 41916
rect 21084 38994 21140 39004
rect 21196 39676 21476 39732
rect 20972 38210 21028 38220
rect 20412 37604 20468 37614
rect 20412 37490 20468 37548
rect 20412 37438 20414 37490
rect 20466 37438 20468 37490
rect 20412 37268 20468 37438
rect 20412 37202 20468 37212
rect 21196 37378 21252 39676
rect 21308 39506 21364 39518
rect 21308 39454 21310 39506
rect 21362 39454 21364 39506
rect 21308 38612 21364 39454
rect 21420 39506 21476 39676
rect 21532 40514 21588 40526
rect 21532 40462 21534 40514
rect 21586 40462 21588 40514
rect 21532 40292 21588 40462
rect 21532 39620 21588 40236
rect 21532 39554 21588 39564
rect 21644 39844 21700 39854
rect 21644 39618 21700 39788
rect 21644 39566 21646 39618
rect 21698 39566 21700 39618
rect 21644 39554 21700 39566
rect 21420 39454 21422 39506
rect 21474 39454 21476 39506
rect 21420 39442 21476 39454
rect 21420 39060 21476 39070
rect 21420 38948 21476 39004
rect 21420 38892 21700 38948
rect 21420 38834 21476 38892
rect 21420 38782 21422 38834
rect 21474 38782 21476 38834
rect 21420 38770 21476 38782
rect 21308 38546 21364 38556
rect 21532 38722 21588 38734
rect 21532 38670 21534 38722
rect 21586 38670 21588 38722
rect 21196 37326 21198 37378
rect 21250 37326 21252 37378
rect 20300 36978 20356 36988
rect 20524 37044 20580 37054
rect 20188 36430 20190 36482
rect 20242 36430 20244 36482
rect 20188 36418 20244 36430
rect 20076 36306 20132 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20300 35924 20356 35934
rect 19964 35028 20020 35038
rect 19964 34934 20020 34972
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20300 34468 20356 35868
rect 20412 34804 20468 34814
rect 20524 34804 20580 36988
rect 20748 36370 20804 36382
rect 20748 36318 20750 36370
rect 20802 36318 20804 36370
rect 20412 34802 20580 34804
rect 20412 34750 20414 34802
rect 20466 34750 20580 34802
rect 20412 34748 20580 34750
rect 20636 35028 20692 35038
rect 20748 35028 20804 36318
rect 20972 36036 21028 36046
rect 20972 35698 21028 35980
rect 20972 35646 20974 35698
rect 21026 35646 21028 35698
rect 20972 35634 21028 35646
rect 21196 35028 21252 37326
rect 21532 37380 21588 38670
rect 21644 38162 21700 38892
rect 21644 38110 21646 38162
rect 21698 38110 21700 38162
rect 21644 38098 21700 38110
rect 21980 37828 22036 41244
rect 22092 41356 22708 41412
rect 22092 41298 22148 41356
rect 22092 41246 22094 41298
rect 22146 41246 22148 41298
rect 22092 41234 22148 41246
rect 22428 41186 22484 41198
rect 22428 41134 22430 41186
rect 22482 41134 22484 41186
rect 22316 41074 22372 41086
rect 22316 41022 22318 41074
rect 22370 41022 22372 41074
rect 22316 40628 22372 41022
rect 22428 41076 22484 41134
rect 22428 41010 22484 41020
rect 22316 40562 22372 40572
rect 22428 40404 22484 40414
rect 22428 40290 22484 40348
rect 22428 40238 22430 40290
rect 22482 40238 22484 40290
rect 22428 40226 22484 40238
rect 22652 39060 22708 41356
rect 22764 40852 22820 44156
rect 22876 42980 22932 45332
rect 23100 44772 23156 45838
rect 23324 44884 23380 46844
rect 23772 46900 23828 46910
rect 23772 46806 23828 46844
rect 23660 46788 23716 46798
rect 23660 46694 23716 46732
rect 23884 46788 23940 46798
rect 23884 46694 23940 46732
rect 23884 46228 23940 46238
rect 23996 46228 24052 47180
rect 23940 46172 24052 46228
rect 24108 46900 24164 47180
rect 24220 47124 24276 47294
rect 24444 47068 24500 47406
rect 24220 47058 24276 47068
rect 24332 47012 24500 47068
rect 24220 46900 24276 46910
rect 24108 46898 24276 46900
rect 24108 46846 24222 46898
rect 24274 46846 24276 46898
rect 24108 46844 24276 46846
rect 23884 46162 23940 46172
rect 23436 46116 23492 46126
rect 23436 45890 23492 46060
rect 23436 45838 23438 45890
rect 23490 45838 23492 45890
rect 23436 45826 23492 45838
rect 23772 45890 23828 45902
rect 23772 45838 23774 45890
rect 23826 45838 23828 45890
rect 23436 44884 23492 44894
rect 23324 44828 23436 44884
rect 23436 44818 23492 44828
rect 23660 44884 23716 44894
rect 23660 44790 23716 44828
rect 23100 44706 23156 44716
rect 23660 44548 23716 44558
rect 23660 44324 23716 44492
rect 23660 44230 23716 44268
rect 23324 44212 23380 44222
rect 22876 42914 22932 42924
rect 22988 44098 23044 44110
rect 22988 44046 22990 44098
rect 23042 44046 23044 44098
rect 22988 43428 23044 44046
rect 23324 43540 23380 44156
rect 23324 43474 23380 43484
rect 23548 44100 23604 44110
rect 23548 43538 23604 44044
rect 23548 43486 23550 43538
rect 23602 43486 23604 43538
rect 23548 43474 23604 43486
rect 22876 42196 22932 42206
rect 22876 42082 22932 42140
rect 22876 42030 22878 42082
rect 22930 42030 22932 42082
rect 22876 42018 22932 42030
rect 22988 42084 23044 43372
rect 23436 42980 23492 42990
rect 23436 42866 23492 42924
rect 23772 42868 23828 45838
rect 23884 45108 23940 45118
rect 24108 45108 24164 46844
rect 24220 46834 24276 46844
rect 24332 45556 24388 47012
rect 24444 46786 24500 46798
rect 24444 46734 24446 46786
rect 24498 46734 24500 46786
rect 24444 46564 24500 46734
rect 24556 46788 24612 46798
rect 24556 46694 24612 46732
rect 24444 46498 24500 46508
rect 24444 45556 24500 45566
rect 24332 45500 24444 45556
rect 24444 45490 24500 45500
rect 24444 45220 24500 45230
rect 24444 45126 24500 45164
rect 23884 45106 24164 45108
rect 23884 45054 23886 45106
rect 23938 45054 24164 45106
rect 23884 45052 24164 45054
rect 24332 45108 24388 45118
rect 23884 45042 23940 45052
rect 24332 45014 24388 45052
rect 24444 44882 24500 44894
rect 24444 44830 24446 44882
rect 24498 44830 24500 44882
rect 24444 44324 24500 44830
rect 24444 44258 24500 44268
rect 24668 44100 24724 47964
rect 24780 47460 24836 47470
rect 24780 47366 24836 47404
rect 24108 44044 24724 44100
rect 23436 42814 23438 42866
rect 23490 42814 23492 42866
rect 23436 42802 23492 42814
rect 23548 42812 23828 42868
rect 23884 43652 23940 43662
rect 23884 43426 23940 43596
rect 23884 43374 23886 43426
rect 23938 43374 23940 43426
rect 22988 42018 23044 42028
rect 23548 42420 23604 42812
rect 23212 41860 23268 41870
rect 23212 41766 23268 41804
rect 22764 39730 22820 40796
rect 22764 39678 22766 39730
rect 22818 39678 22820 39730
rect 22764 39666 22820 39678
rect 22988 40628 23044 40638
rect 22764 39060 22820 39070
rect 22652 39004 22764 39060
rect 21532 37324 21700 37380
rect 21532 37154 21588 37166
rect 21532 37102 21534 37154
rect 21586 37102 21588 37154
rect 21532 36482 21588 37102
rect 21644 37156 21700 37324
rect 21868 37266 21924 37278
rect 21868 37214 21870 37266
rect 21922 37214 21924 37266
rect 21756 37156 21812 37166
rect 21644 37100 21756 37156
rect 21756 37090 21812 37100
rect 21868 36708 21924 37214
rect 21980 37044 22036 37772
rect 21980 36978 22036 36988
rect 22204 37826 22260 37838
rect 22204 37774 22206 37826
rect 22258 37774 22260 37826
rect 21868 36642 21924 36652
rect 21532 36430 21534 36482
rect 21586 36430 21588 36482
rect 21532 36418 21588 36430
rect 21756 36484 21812 36494
rect 21420 35698 21476 35710
rect 21420 35646 21422 35698
rect 21474 35646 21476 35698
rect 21420 35588 21476 35646
rect 21420 35522 21476 35532
rect 21756 35474 21812 36428
rect 21756 35422 21758 35474
rect 21810 35422 21812 35474
rect 21756 35410 21812 35422
rect 21868 35586 21924 35598
rect 21868 35534 21870 35586
rect 21922 35534 21924 35586
rect 21868 35476 21924 35534
rect 21868 35410 21924 35420
rect 21756 35028 21812 35038
rect 20748 35026 21812 35028
rect 20748 34974 21758 35026
rect 21810 34974 21812 35026
rect 20748 34972 21812 34974
rect 20412 34738 20468 34748
rect 20300 34402 20356 34412
rect 19852 34244 19908 34254
rect 19852 34150 19908 34188
rect 19292 33964 19684 34020
rect 20188 34130 20244 34142
rect 20188 34078 20190 34130
rect 20242 34078 20244 34130
rect 19292 33458 19348 33964
rect 19516 33572 19572 33610
rect 19516 33506 19572 33516
rect 19292 33406 19294 33458
rect 19346 33406 19348 33458
rect 19292 33394 19348 33406
rect 19068 32622 19070 32674
rect 19122 32622 19124 32674
rect 18732 32508 19012 32564
rect 17948 32398 17950 32450
rect 18002 32398 18004 32450
rect 17948 32386 18004 32398
rect 16716 31220 16772 31230
rect 16716 31106 16772 31164
rect 16716 31054 16718 31106
rect 16770 31054 16772 31106
rect 16716 31042 16772 31054
rect 16604 30382 16606 30434
rect 16658 30382 16660 30434
rect 16604 30370 16660 30382
rect 15820 30158 15822 30210
rect 15874 30158 15876 30210
rect 15820 30146 15876 30158
rect 16492 30210 16548 30222
rect 16492 30158 16494 30210
rect 16546 30158 16548 30210
rect 15260 29894 15316 29932
rect 16492 29988 16548 30158
rect 17164 30212 17220 31836
rect 18284 31892 18340 31902
rect 18284 31218 18340 31836
rect 18844 31892 18900 31902
rect 18844 31798 18900 31836
rect 18956 31220 19012 32508
rect 19068 31892 19124 32622
rect 19068 31826 19124 31836
rect 19180 33236 19236 33246
rect 18284 31166 18286 31218
rect 18338 31166 18340 31218
rect 18284 31154 18340 31166
rect 18620 31218 19012 31220
rect 18620 31166 18958 31218
rect 19010 31166 19012 31218
rect 18620 31164 19012 31166
rect 18060 31108 18116 31118
rect 18060 30996 18116 31052
rect 17724 30994 18116 30996
rect 17724 30942 18062 30994
rect 18114 30942 18116 30994
rect 17724 30940 18116 30942
rect 17388 30324 17444 30334
rect 17388 30212 17444 30268
rect 17164 30210 17444 30212
rect 17164 30158 17390 30210
rect 17442 30158 17444 30210
rect 17164 30156 17444 30158
rect 17388 30146 17444 30156
rect 16492 28868 16548 29932
rect 17724 30098 17780 30940
rect 18060 30930 18116 30940
rect 18172 30996 18228 31006
rect 18172 30902 18228 30940
rect 17948 30324 18004 30334
rect 17836 30212 17892 30222
rect 17836 30118 17892 30156
rect 17948 30210 18004 30268
rect 17948 30158 17950 30210
rect 18002 30158 18004 30210
rect 17948 30146 18004 30158
rect 18620 30210 18676 31164
rect 18956 31154 19012 31164
rect 19180 31220 19236 33180
rect 20188 33236 20244 34078
rect 20636 34132 20692 34972
rect 21756 34962 21812 34972
rect 22204 34916 22260 37774
rect 22652 35308 22708 39004
rect 22764 38966 22820 39004
rect 22988 38834 23044 40572
rect 23212 39396 23268 39406
rect 23212 39302 23268 39340
rect 22988 38782 22990 38834
rect 23042 38782 23044 38834
rect 22988 38770 23044 38782
rect 23436 38836 23492 38846
rect 23212 38722 23268 38734
rect 23212 38670 23214 38722
rect 23266 38670 23268 38722
rect 22876 38164 22932 38174
rect 22876 38070 22932 38108
rect 22764 38052 22820 38062
rect 22764 37716 22820 37996
rect 23212 38052 23268 38670
rect 23212 37986 23268 37996
rect 23324 38164 23380 38174
rect 23212 37828 23268 37838
rect 23324 37828 23380 38108
rect 23212 37826 23380 37828
rect 23212 37774 23214 37826
rect 23266 37774 23380 37826
rect 23212 37772 23380 37774
rect 23212 37762 23268 37772
rect 22764 37266 22820 37660
rect 22764 37214 22766 37266
rect 22818 37214 22820 37266
rect 22764 37202 22820 37214
rect 22764 37044 22820 37054
rect 22764 36482 22820 36988
rect 22764 36430 22766 36482
rect 22818 36430 22820 36482
rect 22764 36418 22820 36430
rect 22204 34850 22260 34860
rect 22540 35252 22708 35308
rect 23212 35698 23268 35710
rect 23212 35646 23214 35698
rect 23266 35646 23268 35698
rect 22540 35028 22596 35252
rect 20300 33572 20356 33582
rect 20300 33458 20356 33516
rect 20300 33406 20302 33458
rect 20354 33406 20356 33458
rect 20300 33348 20356 33406
rect 20300 33282 20356 33292
rect 20188 33170 20244 33180
rect 19292 33124 19348 33134
rect 19292 33030 19348 33068
rect 19836 32956 20100 32966
rect 19404 32900 19460 32910
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19292 32788 19348 32798
rect 19292 31780 19348 32732
rect 19404 32562 19460 32844
rect 20636 32788 20692 34076
rect 20748 34690 20804 34702
rect 20748 34638 20750 34690
rect 20802 34638 20804 34690
rect 20748 33348 20804 34638
rect 21308 34690 21364 34702
rect 21308 34638 21310 34690
rect 21362 34638 21364 34690
rect 20972 34020 21028 34030
rect 20972 33926 21028 33964
rect 21308 33572 21364 34638
rect 22316 34690 22372 34702
rect 22316 34638 22318 34690
rect 22370 34638 22372 34690
rect 22316 34244 22372 34638
rect 21756 33684 21812 33694
rect 21756 33572 21812 33628
rect 22316 33684 22372 34188
rect 22316 33618 22372 33628
rect 21756 33516 21924 33572
rect 21308 33506 21364 33516
rect 21756 33348 21812 33358
rect 20748 33282 20804 33292
rect 21644 33292 21756 33348
rect 20748 33124 20804 33134
rect 20748 33030 20804 33068
rect 20748 32788 20804 32798
rect 21532 32788 21588 32798
rect 20636 32786 21476 32788
rect 20636 32734 20750 32786
rect 20802 32734 21476 32786
rect 20636 32732 21476 32734
rect 20748 32722 20804 32732
rect 19404 32510 19406 32562
rect 19458 32510 19460 32562
rect 19404 32498 19460 32510
rect 19964 32564 20020 32574
rect 19964 32470 20020 32508
rect 21308 32564 21364 32574
rect 19292 31714 19348 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 18732 30994 18788 31006
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18732 30772 18788 30942
rect 19180 30994 19236 31164
rect 19740 31220 19796 31230
rect 19740 31126 19796 31164
rect 20300 31220 20356 31230
rect 20300 31126 20356 31164
rect 19628 31108 19684 31118
rect 19628 31014 19684 31052
rect 19180 30942 19182 30994
rect 19234 30942 19236 30994
rect 19180 30930 19236 30942
rect 21308 30994 21364 32508
rect 21420 32562 21476 32732
rect 21420 32510 21422 32562
rect 21474 32510 21476 32562
rect 21420 32498 21476 32510
rect 21532 32450 21588 32732
rect 21644 32562 21700 33292
rect 21756 33282 21812 33292
rect 21756 33124 21812 33134
rect 21868 33124 21924 33516
rect 21756 33122 21924 33124
rect 21756 33070 21758 33122
rect 21810 33070 21924 33122
rect 21756 33068 21924 33070
rect 22092 33346 22148 33358
rect 22092 33294 22094 33346
rect 22146 33294 22148 33346
rect 21756 33058 21812 33068
rect 21644 32510 21646 32562
rect 21698 32510 21700 32562
rect 21644 32498 21700 32510
rect 21532 32398 21534 32450
rect 21586 32398 21588 32450
rect 21532 31668 21588 32398
rect 22092 32340 22148 33294
rect 21868 32284 22148 32340
rect 22204 33124 22260 33134
rect 21756 32116 21812 32126
rect 21868 32116 21924 32284
rect 21812 32060 21924 32116
rect 21756 31890 21812 32060
rect 21756 31838 21758 31890
rect 21810 31838 21812 31890
rect 21756 31826 21812 31838
rect 21980 31668 22036 31678
rect 21532 31666 22036 31668
rect 21532 31614 21982 31666
rect 22034 31614 22036 31666
rect 21532 31612 22036 31614
rect 21980 31602 22036 31612
rect 22204 31218 22260 33068
rect 22428 32788 22484 32798
rect 22428 32694 22484 32732
rect 22540 31890 22596 34972
rect 22764 34802 22820 34814
rect 22764 34750 22766 34802
rect 22818 34750 22820 34802
rect 22652 34132 22708 34142
rect 22764 34132 22820 34750
rect 23212 34356 23268 35646
rect 23436 35700 23492 38780
rect 23548 38668 23604 42364
rect 23660 42644 23716 42654
rect 23660 42084 23716 42588
rect 23660 42018 23716 42028
rect 23772 42530 23828 42542
rect 23772 42478 23774 42530
rect 23826 42478 23828 42530
rect 23772 41748 23828 42478
rect 23772 41682 23828 41692
rect 23884 41300 23940 43374
rect 23996 42530 24052 42542
rect 23996 42478 23998 42530
rect 24050 42478 24052 42530
rect 23996 41412 24052 42478
rect 23996 41346 24052 41356
rect 23660 41244 23940 41300
rect 23660 39172 23716 41244
rect 24108 41188 24164 44044
rect 24892 43540 24948 50372
rect 25116 48132 25172 51326
rect 25228 50932 25284 51548
rect 25228 50594 25284 50876
rect 25340 51380 25396 51390
rect 25340 50818 25396 51324
rect 25452 50932 25508 53566
rect 25900 53508 25956 53518
rect 25900 53414 25956 53452
rect 25564 52500 25620 52510
rect 25564 52162 25620 52444
rect 25564 52110 25566 52162
rect 25618 52110 25620 52162
rect 25564 52098 25620 52110
rect 25676 51604 25732 51614
rect 25676 51510 25732 51548
rect 25564 51378 25620 51390
rect 25564 51326 25566 51378
rect 25618 51326 25620 51378
rect 25564 51156 25620 51326
rect 25788 51380 25844 51390
rect 25788 51286 25844 51324
rect 25564 51090 25620 51100
rect 25452 50876 25844 50932
rect 25340 50766 25342 50818
rect 25394 50766 25396 50818
rect 25340 50754 25396 50766
rect 25228 50542 25230 50594
rect 25282 50542 25284 50594
rect 25228 50530 25284 50542
rect 25564 50596 25620 50634
rect 25564 50530 25620 50540
rect 25340 49922 25396 49934
rect 25340 49870 25342 49922
rect 25394 49870 25396 49922
rect 25228 49810 25284 49822
rect 25228 49758 25230 49810
rect 25282 49758 25284 49810
rect 25228 49700 25284 49758
rect 25228 49634 25284 49644
rect 25228 49476 25284 49486
rect 25340 49476 25396 49870
rect 25284 49420 25396 49476
rect 25452 49698 25508 49710
rect 25452 49646 25454 49698
rect 25506 49646 25508 49698
rect 25228 49410 25284 49420
rect 25452 49026 25508 49646
rect 25452 48974 25454 49026
rect 25506 48974 25508 49026
rect 25452 48962 25508 48974
rect 25788 48466 25844 50876
rect 25788 48414 25790 48466
rect 25842 48414 25844 48466
rect 25788 48402 25844 48414
rect 25900 48354 25956 48366
rect 25900 48302 25902 48354
rect 25954 48302 25956 48354
rect 25900 48244 25956 48302
rect 25900 48178 25956 48188
rect 25116 48066 25172 48076
rect 25340 48130 25396 48142
rect 25340 48078 25342 48130
rect 25394 48078 25396 48130
rect 25340 47682 25396 48078
rect 25340 47630 25342 47682
rect 25394 47630 25396 47682
rect 25340 47618 25396 47630
rect 25564 48132 25620 48142
rect 25228 47348 25284 47358
rect 25004 47124 25060 47134
rect 25004 45332 25060 47068
rect 25228 46900 25284 47292
rect 25340 47236 25396 47246
rect 25340 47234 25508 47236
rect 25340 47182 25342 47234
rect 25394 47182 25508 47234
rect 25340 47180 25508 47182
rect 25340 47170 25396 47180
rect 25340 46900 25396 46910
rect 25228 46844 25340 46900
rect 25340 46806 25396 46844
rect 25228 45780 25284 45790
rect 25228 45686 25284 45724
rect 25340 45332 25396 45342
rect 25004 45276 25172 45332
rect 25004 44884 25060 44894
rect 25004 44322 25060 44828
rect 25004 44270 25006 44322
rect 25058 44270 25060 44322
rect 25004 44258 25060 44270
rect 25116 44100 25172 45276
rect 25340 45218 25396 45276
rect 25340 45166 25342 45218
rect 25394 45166 25396 45218
rect 25340 45154 25396 45166
rect 25452 44884 25508 47180
rect 25452 44818 25508 44828
rect 25340 44324 25396 44334
rect 25340 44230 25396 44268
rect 24332 43484 24948 43540
rect 25004 44044 25172 44100
rect 24220 42756 24276 42766
rect 24220 42642 24276 42700
rect 24220 42590 24222 42642
rect 24274 42590 24276 42642
rect 24220 42578 24276 42590
rect 24332 42308 24388 43484
rect 25004 43428 25060 44044
rect 25564 43652 25620 48076
rect 25676 48020 25732 48030
rect 25676 47926 25732 47964
rect 25676 47684 25732 47694
rect 25676 47234 25732 47628
rect 25676 47182 25678 47234
rect 25730 47182 25732 47234
rect 25676 45892 25732 47182
rect 26012 47236 26068 54796
rect 26348 54626 26404 55020
rect 26348 54574 26350 54626
rect 26402 54574 26404 54626
rect 26348 54562 26404 54574
rect 26124 53732 26180 53742
rect 26460 53732 26516 55134
rect 26124 53730 26516 53732
rect 26124 53678 26126 53730
rect 26178 53678 26516 53730
rect 26124 53676 26516 53678
rect 26572 55076 26628 55086
rect 26684 55076 26740 55412
rect 29372 55410 29540 55412
rect 29372 55358 29374 55410
rect 29426 55358 29540 55410
rect 29372 55356 29540 55358
rect 29372 55346 29428 55356
rect 27804 55186 27860 55198
rect 27804 55134 27806 55186
rect 27858 55134 27860 55186
rect 26572 55074 26740 55076
rect 26572 55022 26574 55074
rect 26626 55022 26740 55074
rect 26572 55020 26740 55022
rect 26796 55074 26852 55086
rect 26796 55022 26798 55074
rect 26850 55022 26852 55074
rect 26124 53666 26180 53676
rect 26572 53620 26628 55020
rect 26796 54514 26852 55022
rect 27468 55076 27524 55086
rect 27804 55076 27860 55134
rect 27524 55020 27860 55076
rect 27916 55076 27972 55086
rect 27468 54982 27524 55020
rect 27916 54982 27972 55020
rect 28028 55074 28084 55086
rect 28028 55022 28030 55074
rect 28082 55022 28084 55074
rect 27244 54738 27300 54750
rect 27244 54686 27246 54738
rect 27298 54686 27300 54738
rect 26796 54462 26798 54514
rect 26850 54462 26852 54514
rect 26796 54450 26852 54462
rect 27132 54516 27188 54526
rect 27132 54422 27188 54460
rect 27244 54292 27300 54686
rect 28028 54740 28084 55022
rect 28588 55074 28644 55086
rect 28588 55022 28590 55074
rect 28642 55022 28644 55074
rect 28588 54852 28644 55022
rect 28588 54786 28644 54796
rect 29372 54852 29428 54862
rect 28028 54516 28084 54684
rect 29372 54626 29428 54796
rect 29372 54574 29374 54626
rect 29426 54574 29428 54626
rect 28140 54516 28196 54526
rect 28028 54514 28196 54516
rect 28028 54462 28142 54514
rect 28194 54462 28196 54514
rect 28028 54460 28196 54462
rect 27916 54404 27972 54414
rect 27244 54226 27300 54236
rect 27804 54402 27972 54404
rect 27804 54350 27918 54402
rect 27970 54350 27972 54402
rect 27804 54348 27972 54350
rect 27804 54068 27860 54348
rect 27916 54338 27972 54348
rect 26348 53564 26628 53620
rect 27020 53618 27076 53630
rect 27020 53566 27022 53618
rect 27074 53566 27076 53618
rect 26124 49810 26180 49822
rect 26124 49758 26126 49810
rect 26178 49758 26180 49810
rect 26124 48580 26180 49758
rect 26124 47460 26180 48524
rect 26124 47394 26180 47404
rect 26236 49026 26292 49038
rect 26236 48974 26238 49026
rect 26290 48974 26292 49026
rect 26124 47236 26180 47246
rect 26012 47234 26180 47236
rect 26012 47182 26126 47234
rect 26178 47182 26180 47234
rect 26012 47180 26180 47182
rect 25900 46900 25956 46910
rect 25788 46562 25844 46574
rect 25788 46510 25790 46562
rect 25842 46510 25844 46562
rect 25788 46452 25844 46510
rect 25788 46386 25844 46396
rect 25676 45826 25732 45836
rect 25788 45444 25844 45454
rect 25676 45106 25732 45118
rect 25676 45054 25678 45106
rect 25730 45054 25732 45106
rect 25676 44884 25732 45054
rect 25676 44818 25732 44828
rect 25564 43596 25732 43652
rect 25228 43540 25284 43550
rect 25228 43446 25284 43484
rect 24444 43372 25060 43428
rect 25564 43428 25620 43438
rect 24444 42532 24500 43372
rect 25564 43334 25620 43372
rect 25452 43316 25508 43326
rect 25452 43222 25508 43260
rect 24556 42924 25172 42980
rect 24556 42866 24612 42924
rect 24556 42814 24558 42866
rect 24610 42814 24612 42866
rect 24556 42802 24612 42814
rect 24668 42756 24724 42766
rect 24668 42662 24724 42700
rect 24892 42756 24948 42766
rect 24444 42530 24612 42532
rect 24444 42478 24446 42530
rect 24498 42478 24612 42530
rect 24444 42476 24612 42478
rect 24444 42466 24500 42476
rect 24556 42308 24612 42476
rect 24332 42252 24500 42308
rect 23660 39106 23716 39116
rect 23772 41132 24164 41188
rect 24220 41970 24276 41982
rect 24220 41918 24222 41970
rect 24274 41918 24276 41970
rect 23660 38836 23716 38846
rect 23660 38742 23716 38780
rect 23548 38612 23716 38668
rect 23548 37828 23604 37838
rect 23548 37734 23604 37772
rect 23548 36484 23604 36494
rect 23548 36390 23604 36428
rect 23660 36036 23716 38612
rect 23772 38052 23828 41132
rect 24108 40516 24164 40526
rect 24108 40402 24164 40460
rect 24108 40350 24110 40402
rect 24162 40350 24164 40402
rect 24108 40338 24164 40350
rect 24108 39732 24164 39742
rect 24108 39638 24164 39676
rect 23884 39618 23940 39630
rect 23884 39566 23886 39618
rect 23938 39566 23940 39618
rect 23884 38274 23940 39566
rect 24220 39620 24276 41918
rect 24220 39618 24388 39620
rect 24220 39566 24222 39618
rect 24274 39566 24388 39618
rect 24220 39564 24388 39566
rect 24220 39554 24276 39564
rect 24220 39396 24276 39406
rect 23996 39060 24052 39070
rect 23996 38834 24052 39004
rect 24108 38948 24164 38958
rect 24108 38854 24164 38892
rect 23996 38782 23998 38834
rect 24050 38782 24052 38834
rect 23996 38770 24052 38782
rect 23884 38222 23886 38274
rect 23938 38222 23940 38274
rect 23884 38210 23940 38222
rect 24108 38164 24164 38174
rect 23772 37996 23940 38052
rect 23772 37826 23828 37838
rect 23772 37774 23774 37826
rect 23826 37774 23828 37826
rect 23772 37492 23828 37774
rect 23772 37426 23828 37436
rect 23660 35970 23716 35980
rect 23548 35924 23604 35934
rect 23548 35830 23604 35868
rect 23436 35634 23492 35644
rect 23436 34916 23492 34926
rect 23548 34916 23604 34926
rect 23492 34914 23604 34916
rect 23492 34862 23550 34914
rect 23602 34862 23604 34914
rect 23492 34860 23604 34862
rect 23212 34300 23380 34356
rect 23212 34132 23268 34142
rect 22764 34130 23268 34132
rect 22764 34078 23214 34130
rect 23266 34078 23268 34130
rect 22764 34076 23268 34078
rect 22652 34038 22708 34076
rect 23212 33908 23268 34076
rect 23212 33842 23268 33852
rect 22876 33796 22932 33806
rect 22652 33348 22708 33358
rect 22652 33254 22708 33292
rect 22876 32676 22932 33740
rect 23212 33458 23268 33470
rect 23212 33406 23214 33458
rect 23266 33406 23268 33458
rect 22876 32582 22932 32620
rect 23100 33348 23156 33358
rect 22540 31838 22542 31890
rect 22594 31838 22596 31890
rect 22540 31826 22596 31838
rect 23100 31668 23156 33292
rect 23212 33012 23268 33406
rect 23324 33348 23380 34300
rect 23324 33282 23380 33292
rect 23436 33684 23492 34860
rect 23548 34850 23604 34860
rect 23772 34244 23828 34254
rect 23884 34244 23940 37996
rect 24108 38050 24164 38108
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 24108 37940 24164 37998
rect 24108 35588 24164 37884
rect 24220 37268 24276 39340
rect 24332 38388 24388 39564
rect 24332 38322 24388 38332
rect 24444 38612 24500 42252
rect 24556 42242 24612 42252
rect 24780 41972 24836 41982
rect 24668 41916 24780 41972
rect 24556 41748 24612 41758
rect 24556 41654 24612 41692
rect 24668 41186 24724 41916
rect 24780 41878 24836 41916
rect 24892 41298 24948 42700
rect 24892 41246 24894 41298
rect 24946 41246 24948 41298
rect 24892 41234 24948 41246
rect 24668 41134 24670 41186
rect 24722 41134 24724 41186
rect 24668 41122 24724 41134
rect 25004 41186 25060 41198
rect 25004 41134 25006 41186
rect 25058 41134 25060 41186
rect 24444 38164 24500 38556
rect 24444 38098 24500 38108
rect 24556 40516 24612 40526
rect 24332 37938 24388 37950
rect 24332 37886 24334 37938
rect 24386 37886 24388 37938
rect 24332 37828 24388 37886
rect 24332 37604 24388 37772
rect 24332 37538 24388 37548
rect 24444 37826 24500 37838
rect 24444 37774 24446 37826
rect 24498 37774 24500 37826
rect 24332 37268 24388 37278
rect 24220 37212 24332 37268
rect 24332 37174 24388 37212
rect 24444 36932 24500 37774
rect 24444 36866 24500 36876
rect 24556 36708 24612 40460
rect 24668 40404 24724 40414
rect 25004 40404 25060 41134
rect 24668 40402 25060 40404
rect 24668 40350 24670 40402
rect 24722 40350 25060 40402
rect 24668 40348 25060 40350
rect 24668 40338 24724 40348
rect 24668 38724 24724 38762
rect 24668 38658 24724 38668
rect 24668 37828 24724 37838
rect 24668 37734 24724 37772
rect 24780 37716 24836 40348
rect 24892 39508 24948 39518
rect 24892 39414 24948 39452
rect 25004 38164 25060 38174
rect 25004 38070 25060 38108
rect 24892 38052 24948 38062
rect 24892 37958 24948 37996
rect 25116 38050 25172 42924
rect 25676 42644 25732 43596
rect 25788 42866 25844 45388
rect 25788 42814 25790 42866
rect 25842 42814 25844 42866
rect 25788 42802 25844 42814
rect 25676 42578 25732 42588
rect 25228 42530 25284 42542
rect 25228 42478 25230 42530
rect 25282 42478 25284 42530
rect 25228 42420 25284 42478
rect 25228 42354 25284 42364
rect 25564 42308 25620 42318
rect 25452 42084 25508 42094
rect 25228 41412 25284 41422
rect 25228 40402 25284 41356
rect 25340 40516 25396 40526
rect 25340 40422 25396 40460
rect 25228 40350 25230 40402
rect 25282 40350 25284 40402
rect 25228 40338 25284 40350
rect 25452 40292 25508 42028
rect 25340 40236 25508 40292
rect 25564 41858 25620 42252
rect 25900 42196 25956 46844
rect 26124 45332 26180 47180
rect 26124 45266 26180 45276
rect 26012 45218 26068 45230
rect 26012 45166 26014 45218
rect 26066 45166 26068 45218
rect 26012 44324 26068 45166
rect 26236 45108 26292 48974
rect 26348 47908 26404 53564
rect 26908 53508 26964 53518
rect 26908 53414 26964 53452
rect 26796 53284 26852 53294
rect 26460 52834 26516 52846
rect 26460 52782 26462 52834
rect 26514 52782 26516 52834
rect 26460 52500 26516 52782
rect 26460 52434 26516 52444
rect 26460 51380 26516 51390
rect 26516 51324 26628 51380
rect 26460 51286 26516 51324
rect 26460 50484 26516 50494
rect 26460 50390 26516 50428
rect 26572 49364 26628 51324
rect 26684 49810 26740 49822
rect 26684 49758 26686 49810
rect 26738 49758 26740 49810
rect 26684 49700 26740 49758
rect 26684 49634 26740 49644
rect 26572 49308 26740 49364
rect 26460 48914 26516 48926
rect 26460 48862 26462 48914
rect 26514 48862 26516 48914
rect 26460 48468 26516 48862
rect 26460 48402 26516 48412
rect 26460 48244 26516 48254
rect 26460 48150 26516 48188
rect 26348 47842 26404 47852
rect 26684 47460 26740 49308
rect 26236 45042 26292 45052
rect 26348 47404 26740 47460
rect 26796 47682 26852 53228
rect 26908 52164 26964 52174
rect 26908 52070 26964 52108
rect 26908 51266 26964 51278
rect 26908 51214 26910 51266
rect 26962 51214 26964 51266
rect 26908 50484 26964 51214
rect 26908 49476 26964 50428
rect 26908 49410 26964 49420
rect 27020 50034 27076 53566
rect 27692 53508 27748 53518
rect 27580 53452 27692 53508
rect 27356 52276 27412 52286
rect 27020 49982 27022 50034
rect 27074 49982 27076 50034
rect 27020 49028 27076 49982
rect 27132 52050 27188 52062
rect 27132 51998 27134 52050
rect 27186 51998 27188 52050
rect 27132 49924 27188 51998
rect 27244 51940 27300 51950
rect 27244 51846 27300 51884
rect 27132 49252 27188 49868
rect 27132 49186 27188 49196
rect 27244 51378 27300 51390
rect 27244 51326 27246 51378
rect 27298 51326 27300 51378
rect 27244 51156 27300 51326
rect 27020 48962 27076 48972
rect 27132 48802 27188 48814
rect 27132 48750 27134 48802
rect 27186 48750 27188 48802
rect 27132 48468 27188 48750
rect 27132 48402 27188 48412
rect 27244 48354 27300 51100
rect 27356 50596 27412 52220
rect 27356 50530 27412 50540
rect 27468 52274 27524 52286
rect 27468 52222 27470 52274
rect 27522 52222 27524 52274
rect 27468 50484 27524 52222
rect 27580 51828 27636 53452
rect 27692 53414 27748 53452
rect 27804 53170 27860 54012
rect 27916 53732 27972 53742
rect 28028 53732 28084 54460
rect 28140 54450 28196 54460
rect 28476 54516 28532 54526
rect 29036 54516 29092 54526
rect 28476 54514 29092 54516
rect 28476 54462 28478 54514
rect 28530 54462 29038 54514
rect 29090 54462 29092 54514
rect 28476 54460 29092 54462
rect 28476 54450 28532 54460
rect 28476 53844 28532 53854
rect 28476 53750 28532 53788
rect 27916 53730 28084 53732
rect 27916 53678 27918 53730
rect 27970 53678 28084 53730
rect 27916 53676 28084 53678
rect 27916 53666 27972 53676
rect 28364 53618 28420 53630
rect 28364 53566 28366 53618
rect 28418 53566 28420 53618
rect 28140 53506 28196 53518
rect 28140 53454 28142 53506
rect 28194 53454 28196 53506
rect 28140 53284 28196 53454
rect 28252 53508 28308 53518
rect 28364 53508 28420 53566
rect 29036 53620 29092 54460
rect 29372 53730 29428 54574
rect 29372 53678 29374 53730
rect 29426 53678 29428 53730
rect 29260 53620 29316 53630
rect 29036 53618 29316 53620
rect 29036 53566 29262 53618
rect 29314 53566 29316 53618
rect 29036 53564 29316 53566
rect 29260 53554 29316 53564
rect 28308 53452 28420 53508
rect 28252 53442 28308 53452
rect 28140 53218 28196 53228
rect 28812 53284 28868 53294
rect 27804 53118 27806 53170
rect 27858 53118 27860 53170
rect 27804 53106 27860 53118
rect 28812 53170 28868 53228
rect 28812 53118 28814 53170
rect 28866 53118 28868 53170
rect 28812 53106 28868 53118
rect 28140 53060 28196 53070
rect 28588 53060 28644 53070
rect 28140 53058 28308 53060
rect 28140 53006 28142 53058
rect 28194 53006 28308 53058
rect 28140 53004 28308 53006
rect 28140 52994 28196 53004
rect 27692 52162 27748 52174
rect 27692 52110 27694 52162
rect 27746 52110 27748 52162
rect 27692 52052 27748 52110
rect 27692 51986 27748 51996
rect 27580 51772 27748 51828
rect 27692 51044 27748 51772
rect 28252 51492 28308 53004
rect 28252 51426 28308 51436
rect 28364 52050 28420 52062
rect 28364 51998 28366 52050
rect 28418 51998 28420 52050
rect 28364 51490 28420 51998
rect 28364 51438 28366 51490
rect 28418 51438 28420 51490
rect 27804 51380 27860 51390
rect 28140 51380 28196 51390
rect 27804 51378 28196 51380
rect 27804 51326 27806 51378
rect 27858 51326 28142 51378
rect 28194 51326 28196 51378
rect 27804 51324 28196 51326
rect 27804 51314 27860 51324
rect 28140 51314 28196 51324
rect 28364 51380 28420 51438
rect 28364 51314 28420 51324
rect 28476 51490 28532 51502
rect 28476 51438 28478 51490
rect 28530 51438 28532 51490
rect 28252 51266 28308 51278
rect 28252 51214 28254 51266
rect 28306 51214 28308 51266
rect 27692 50988 27972 51044
rect 27580 50708 27636 50718
rect 27580 50614 27636 50652
rect 27804 50596 27860 50606
rect 27692 50484 27748 50494
rect 27468 50482 27748 50484
rect 27468 50430 27694 50482
rect 27746 50430 27748 50482
rect 27468 50428 27748 50430
rect 27692 50418 27748 50428
rect 27356 50372 27412 50382
rect 27356 49026 27412 50316
rect 27356 48974 27358 49026
rect 27410 48974 27412 49026
rect 27356 48692 27412 48974
rect 27356 48626 27412 48636
rect 27468 49028 27524 49038
rect 27244 48302 27246 48354
rect 27298 48302 27300 48354
rect 27244 48290 27300 48302
rect 27468 48242 27524 48972
rect 27468 48190 27470 48242
rect 27522 48190 27524 48242
rect 26908 48132 26964 48142
rect 26908 48038 26964 48076
rect 26796 47630 26798 47682
rect 26850 47630 26852 47682
rect 26012 44258 26068 44268
rect 26348 43540 26404 47404
rect 26684 47234 26740 47246
rect 26684 47182 26686 47234
rect 26738 47182 26740 47234
rect 26684 47124 26740 47182
rect 26684 47058 26740 47068
rect 26796 46788 26852 47630
rect 27356 47572 27412 47582
rect 27356 47478 27412 47516
rect 26684 46562 26740 46574
rect 26684 46510 26686 46562
rect 26738 46510 26740 46562
rect 26460 46452 26516 46462
rect 26460 45330 26516 46396
rect 26460 45278 26462 45330
rect 26514 45278 26516 45330
rect 26460 45266 26516 45278
rect 26572 46340 26628 46350
rect 26572 45444 26628 46284
rect 26684 46116 26740 46510
rect 26796 46452 26852 46732
rect 26796 46386 26852 46396
rect 27020 47458 27076 47470
rect 27020 47406 27022 47458
rect 27074 47406 27076 47458
rect 27020 46676 27076 47406
rect 27468 47458 27524 48190
rect 27468 47406 27470 47458
rect 27522 47406 27524 47458
rect 27244 47346 27300 47358
rect 27244 47294 27246 47346
rect 27298 47294 27300 47346
rect 27244 47068 27300 47294
rect 27468 47348 27524 47406
rect 27468 47282 27524 47292
rect 27580 48468 27636 48478
rect 27580 48244 27636 48412
rect 27580 47458 27636 48188
rect 27580 47406 27582 47458
rect 27634 47406 27636 47458
rect 27020 46450 27076 46620
rect 27020 46398 27022 46450
rect 27074 46398 27076 46450
rect 27020 46386 27076 46398
rect 27132 47012 27300 47068
rect 27356 47236 27412 47246
rect 26684 45890 26740 46060
rect 26684 45838 26686 45890
rect 26738 45838 26740 45890
rect 26684 45826 26740 45838
rect 27020 45892 27076 45902
rect 26684 45668 26740 45678
rect 26684 45666 26852 45668
rect 26684 45614 26686 45666
rect 26738 45614 26852 45666
rect 26684 45612 26852 45614
rect 26684 45602 26740 45612
rect 26572 44322 26628 45388
rect 26572 44270 26574 44322
rect 26626 44270 26628 44322
rect 26572 44258 26628 44270
rect 26684 45332 26740 45342
rect 26348 43474 26404 43484
rect 26684 43316 26740 45276
rect 26796 45220 26852 45612
rect 26796 45164 26964 45220
rect 26796 44996 26852 45006
rect 26796 44902 26852 44940
rect 26908 44660 26964 45164
rect 27020 45106 27076 45836
rect 27132 45220 27188 47012
rect 27244 46676 27300 46686
rect 27244 46582 27300 46620
rect 27132 45154 27188 45164
rect 27244 45666 27300 45678
rect 27244 45614 27246 45666
rect 27298 45614 27300 45666
rect 27020 45054 27022 45106
rect 27074 45054 27076 45106
rect 27020 45042 27076 45054
rect 26908 44594 26964 44604
rect 27132 44210 27188 44222
rect 27132 44158 27134 44210
rect 27186 44158 27188 44210
rect 26908 44098 26964 44110
rect 26908 44046 26910 44098
rect 26962 44046 26964 44098
rect 26908 43652 26964 44046
rect 26908 43586 26964 43596
rect 26348 43260 26684 43316
rect 26124 42532 26180 42542
rect 25564 41806 25566 41858
rect 25618 41806 25620 41858
rect 25340 39730 25396 40236
rect 25564 40180 25620 41806
rect 25340 39678 25342 39730
rect 25394 39678 25396 39730
rect 25340 39666 25396 39678
rect 25452 40124 25620 40180
rect 25676 42140 25956 42196
rect 26012 42420 26068 42430
rect 25228 39508 25284 39518
rect 25452 39508 25508 40124
rect 25228 39506 25508 39508
rect 25228 39454 25230 39506
rect 25282 39454 25508 39506
rect 25228 39452 25508 39454
rect 25564 39620 25620 39630
rect 25676 39620 25732 42140
rect 26012 41972 26068 42364
rect 26124 42194 26180 42476
rect 26124 42142 26126 42194
rect 26178 42142 26180 42194
rect 26124 42130 26180 42142
rect 26348 42194 26404 43260
rect 26684 43250 26740 43260
rect 26796 43538 26852 43550
rect 26796 43486 26798 43538
rect 26850 43486 26852 43538
rect 26572 43092 26628 43102
rect 26572 42866 26628 43036
rect 26572 42814 26574 42866
rect 26626 42814 26628 42866
rect 26572 42802 26628 42814
rect 26348 42142 26350 42194
rect 26402 42142 26404 42194
rect 26012 41878 26068 41916
rect 26348 41860 26404 42142
rect 26572 42084 26628 42094
rect 26572 41970 26628 42028
rect 26572 41918 26574 41970
rect 26626 41918 26628 41970
rect 26572 41906 26628 41918
rect 26796 42084 26852 43486
rect 26908 43316 26964 43326
rect 27132 43316 27188 44158
rect 27244 43650 27300 45614
rect 27356 45444 27412 47180
rect 27468 47124 27524 47134
rect 27468 45890 27524 47068
rect 27468 45838 27470 45890
rect 27522 45838 27524 45890
rect 27468 45826 27524 45838
rect 27580 45780 27636 47406
rect 27692 46674 27748 46686
rect 27692 46622 27694 46674
rect 27746 46622 27748 46674
rect 27692 46564 27748 46622
rect 27692 46004 27748 46508
rect 27804 46228 27860 50540
rect 27916 49700 27972 50988
rect 28252 50708 28308 51214
rect 28252 50642 28308 50652
rect 28140 50484 28196 50494
rect 28140 50390 28196 50428
rect 28476 50484 28532 51438
rect 28476 50418 28532 50428
rect 28588 49924 28644 53004
rect 29260 52836 29316 52846
rect 29372 52836 29428 53678
rect 29260 52834 29428 52836
rect 29260 52782 29262 52834
rect 29314 52782 29428 52834
rect 29260 52780 29428 52782
rect 29484 54628 29540 55356
rect 28700 52164 28756 52174
rect 29260 52164 29316 52780
rect 28700 52162 29316 52164
rect 28700 52110 28702 52162
rect 28754 52110 29316 52162
rect 28700 52108 29316 52110
rect 28700 52098 28756 52108
rect 29260 51940 29316 51950
rect 29484 51940 29540 54572
rect 29708 55298 29764 55310
rect 29708 55246 29710 55298
rect 29762 55246 29764 55298
rect 29708 55076 29764 55246
rect 30156 55188 30212 55198
rect 30156 55076 30212 55132
rect 30828 55188 30884 55198
rect 30828 55094 30884 55132
rect 31500 55188 31556 55198
rect 29708 55074 30212 55076
rect 29708 55022 30158 55074
rect 30210 55022 30212 55074
rect 29708 55020 30212 55022
rect 29708 54516 29764 55020
rect 30156 55010 30212 55020
rect 30492 55074 30548 55086
rect 30492 55022 30494 55074
rect 30546 55022 30548 55074
rect 29708 54450 29764 54460
rect 30156 54404 30212 54414
rect 30156 54310 30212 54348
rect 29148 51938 29540 51940
rect 29148 51886 29262 51938
rect 29314 51886 29540 51938
rect 29148 51884 29540 51886
rect 30044 53956 30100 53966
rect 30044 53730 30100 53900
rect 30044 53678 30046 53730
rect 30098 53678 30100 53730
rect 28924 51380 28980 51390
rect 29148 51380 29204 51884
rect 29260 51874 29316 51884
rect 28924 51378 29204 51380
rect 28924 51326 28926 51378
rect 28978 51326 29204 51378
rect 28924 51324 29204 51326
rect 29260 51492 29316 51502
rect 29260 51378 29316 51436
rect 29260 51326 29262 51378
rect 29314 51326 29316 51378
rect 28924 51314 28980 51324
rect 28700 50372 28756 50382
rect 28812 50372 28868 50382
rect 28700 50370 28812 50372
rect 28700 50318 28702 50370
rect 28754 50318 28812 50370
rect 28700 50316 28812 50318
rect 28700 50306 28756 50316
rect 28588 49868 28756 49924
rect 27916 49634 27972 49644
rect 28028 49812 28084 49822
rect 27916 49252 27972 49262
rect 27916 48020 27972 49196
rect 28028 49028 28084 49756
rect 28588 49700 28644 49710
rect 28588 49606 28644 49644
rect 28028 48962 28084 48972
rect 28028 48802 28084 48814
rect 28028 48750 28030 48802
rect 28082 48750 28084 48802
rect 28028 48244 28084 48750
rect 28588 48804 28644 48814
rect 28700 48804 28756 49868
rect 28812 49140 28868 50316
rect 28812 49074 28868 49084
rect 29036 49700 29092 51324
rect 29148 50596 29204 50606
rect 29260 50596 29316 51326
rect 29820 51268 29876 51278
rect 29820 51266 29988 51268
rect 29820 51214 29822 51266
rect 29874 51214 29988 51266
rect 29820 51212 29988 51214
rect 29820 51202 29876 51212
rect 29484 50596 29540 50606
rect 29260 50594 29540 50596
rect 29260 50542 29486 50594
rect 29538 50542 29540 50594
rect 29260 50540 29540 50542
rect 29148 50502 29204 50540
rect 29484 50530 29540 50540
rect 29596 50370 29652 50382
rect 29596 50318 29598 50370
rect 29650 50318 29652 50370
rect 29596 50036 29652 50318
rect 29708 50372 29764 50382
rect 29708 50278 29764 50316
rect 29820 50036 29876 50046
rect 29596 50034 29876 50036
rect 29596 49982 29822 50034
rect 29874 49982 29876 50034
rect 29596 49980 29876 49982
rect 29820 49970 29876 49980
rect 29596 49810 29652 49822
rect 29932 49812 29988 51212
rect 30044 50596 30100 53678
rect 30268 53620 30324 53630
rect 30268 53618 30436 53620
rect 30268 53566 30270 53618
rect 30322 53566 30436 53618
rect 30268 53564 30436 53566
rect 30268 53554 30324 53564
rect 30380 52724 30436 53564
rect 30380 52658 30436 52668
rect 30156 52612 30212 52622
rect 30156 51380 30212 52556
rect 30156 51314 30212 51324
rect 30492 52162 30548 55022
rect 30604 55076 30660 55086
rect 30604 54514 30660 55020
rect 30604 54462 30606 54514
rect 30658 54462 30660 54514
rect 30604 54450 30660 54462
rect 31164 55074 31220 55086
rect 31164 55022 31166 55074
rect 31218 55022 31220 55074
rect 30940 53844 30996 53854
rect 30940 53730 30996 53788
rect 30940 53678 30942 53730
rect 30994 53678 30996 53730
rect 30940 53666 30996 53678
rect 30828 53172 30884 53182
rect 30828 53078 30884 53116
rect 31052 52946 31108 52958
rect 31052 52894 31054 52946
rect 31106 52894 31108 52946
rect 30940 52836 30996 52846
rect 30940 52742 30996 52780
rect 31052 52724 31108 52894
rect 31164 52724 31220 55022
rect 31500 53506 31556 55132
rect 31500 53454 31502 53506
rect 31554 53454 31556 53506
rect 31500 53442 31556 53454
rect 31052 52668 31164 52724
rect 31164 52658 31220 52668
rect 31276 53058 31332 53070
rect 31276 53006 31278 53058
rect 31330 53006 31332 53058
rect 31276 52386 31332 53006
rect 31276 52334 31278 52386
rect 31330 52334 31332 52386
rect 31276 52322 31332 52334
rect 30492 52110 30494 52162
rect 30546 52110 30548 52162
rect 30492 51380 30548 52110
rect 30828 52052 30884 52062
rect 30828 51940 30884 51996
rect 30716 51938 30884 51940
rect 30716 51886 30830 51938
rect 30882 51886 30884 51938
rect 30716 51884 30884 51886
rect 30604 51380 30660 51390
rect 30492 51378 30660 51380
rect 30492 51326 30606 51378
rect 30658 51326 30660 51378
rect 30492 51324 30660 51326
rect 30044 50530 30100 50540
rect 30380 50482 30436 50494
rect 30380 50430 30382 50482
rect 30434 50430 30436 50482
rect 30268 50372 30324 50382
rect 30380 50372 30436 50430
rect 30324 50316 30436 50372
rect 30268 50306 30324 50316
rect 30380 50036 30436 50316
rect 30492 50372 30548 51324
rect 30604 51314 30660 51324
rect 30716 51268 30772 51884
rect 30828 51874 30884 51884
rect 31164 52050 31220 52062
rect 31164 51998 31166 52050
rect 31218 51998 31220 52050
rect 31164 51716 31220 51998
rect 31276 52052 31332 52062
rect 31276 51958 31332 51996
rect 31220 51660 31444 51716
rect 31164 51650 31220 51660
rect 30940 51492 30996 51502
rect 30828 51380 30884 51390
rect 30828 51286 30884 51324
rect 30716 51202 30772 51212
rect 30492 50306 30548 50316
rect 30604 50036 30660 50046
rect 30380 50034 30660 50036
rect 30380 49982 30606 50034
rect 30658 49982 30660 50034
rect 30380 49980 30660 49982
rect 30604 49970 30660 49980
rect 30044 49924 30100 49962
rect 30044 49858 30100 49868
rect 30268 49812 30324 49822
rect 29596 49758 29598 49810
rect 29650 49758 29652 49810
rect 29260 49700 29316 49710
rect 29596 49700 29652 49758
rect 29820 49756 29988 49812
rect 30156 49756 30268 49812
rect 29036 49698 29652 49700
rect 29036 49646 29262 49698
rect 29314 49646 29652 49698
rect 29036 49644 29652 49646
rect 29708 49700 29764 49710
rect 28644 48748 28756 48804
rect 28588 48710 28644 48748
rect 29036 48692 29092 49644
rect 29260 49634 29316 49644
rect 28812 48636 29092 48692
rect 29148 49476 29204 49486
rect 28028 48178 28084 48188
rect 28140 48242 28196 48254
rect 28140 48190 28142 48242
rect 28194 48190 28196 48242
rect 28140 48020 28196 48190
rect 27916 47964 28196 48020
rect 28364 48244 28420 48254
rect 27916 46340 27972 47964
rect 28140 47460 28196 47470
rect 28140 47366 28196 47404
rect 28252 47348 28308 47358
rect 28252 47254 28308 47292
rect 28028 47234 28084 47246
rect 28028 47182 28030 47234
rect 28082 47182 28084 47234
rect 28028 47012 28084 47182
rect 28364 47124 28420 48188
rect 28364 47058 28420 47068
rect 28476 47234 28532 47246
rect 28476 47182 28478 47234
rect 28530 47182 28532 47234
rect 28028 46946 28084 46956
rect 27916 46274 27972 46284
rect 28140 46562 28196 46574
rect 28140 46510 28142 46562
rect 28194 46510 28196 46562
rect 27804 46162 27860 46172
rect 28028 46228 28084 46238
rect 28140 46228 28196 46510
rect 28084 46172 28196 46228
rect 28028 46162 28084 46172
rect 27692 45938 27748 45948
rect 28364 45892 28420 45902
rect 28364 45798 28420 45836
rect 27692 45780 27748 45790
rect 27580 45778 27748 45780
rect 27580 45726 27694 45778
rect 27746 45726 27748 45778
rect 27580 45724 27748 45726
rect 27692 45714 27748 45724
rect 27804 45780 27860 45790
rect 28028 45780 28084 45790
rect 27804 45778 28084 45780
rect 27804 45726 27806 45778
rect 27858 45726 28030 45778
rect 28082 45726 28084 45778
rect 27804 45724 28084 45726
rect 27804 45714 27860 45724
rect 28028 45714 28084 45724
rect 28140 45668 28196 45678
rect 27356 45388 28084 45444
rect 27468 45108 27524 45118
rect 27804 45108 27860 45118
rect 27468 45014 27524 45052
rect 27692 45106 27860 45108
rect 27692 45054 27806 45106
rect 27858 45054 27860 45106
rect 27692 45052 27860 45054
rect 27244 43598 27246 43650
rect 27298 43598 27300 43650
rect 27244 43586 27300 43598
rect 27468 43650 27524 43662
rect 27468 43598 27470 43650
rect 27522 43598 27524 43650
rect 26908 43314 27188 43316
rect 26908 43262 26910 43314
rect 26962 43262 27188 43314
rect 26908 43260 27188 43262
rect 26908 43250 26964 43260
rect 27468 43204 27524 43598
rect 27580 43540 27636 43550
rect 27580 43316 27636 43484
rect 27580 43250 27636 43260
rect 27132 43148 27524 43204
rect 27132 43092 27188 43148
rect 27692 43092 27748 45052
rect 27804 45042 27860 45052
rect 26012 41186 26068 41198
rect 26012 41134 26014 41186
rect 26066 41134 26068 41186
rect 25564 39618 25732 39620
rect 25564 39566 25566 39618
rect 25618 39566 25732 39618
rect 25564 39564 25732 39566
rect 25788 40068 25844 40078
rect 25788 39618 25844 40012
rect 25788 39566 25790 39618
rect 25842 39566 25844 39618
rect 25228 39396 25284 39452
rect 25228 39330 25284 39340
rect 25340 38722 25396 38734
rect 25340 38670 25342 38722
rect 25394 38670 25396 38722
rect 25340 38612 25396 38670
rect 25340 38546 25396 38556
rect 25564 38276 25620 39564
rect 25788 39554 25844 39566
rect 26012 39060 26068 41134
rect 26124 40852 26180 40862
rect 26124 40402 26180 40796
rect 26236 40740 26292 40750
rect 26236 40626 26292 40684
rect 26236 40574 26238 40626
rect 26290 40574 26292 40626
rect 26236 40562 26292 40574
rect 26124 40350 26126 40402
rect 26178 40350 26180 40402
rect 26124 40338 26180 40350
rect 26348 40180 26404 41804
rect 26460 41858 26516 41870
rect 26460 41806 26462 41858
rect 26514 41806 26516 41858
rect 26460 41748 26516 41806
rect 26684 41860 26740 41870
rect 26684 41748 26740 41804
rect 26460 41692 26740 41748
rect 26796 41636 26852 42028
rect 26124 40124 26404 40180
rect 26460 41580 26852 41636
rect 26908 43036 27188 43092
rect 27356 43036 27748 43092
rect 26124 39506 26180 40124
rect 26124 39454 26126 39506
rect 26178 39454 26180 39506
rect 26124 39442 26180 39454
rect 26348 39618 26404 39630
rect 26348 39566 26350 39618
rect 26402 39566 26404 39618
rect 26012 38994 26068 39004
rect 26236 39172 26292 39182
rect 26124 38948 26180 38958
rect 26124 38724 26180 38892
rect 26236 38836 26292 39116
rect 26348 39060 26404 39566
rect 26348 38994 26404 39004
rect 26348 38836 26404 38846
rect 26236 38834 26404 38836
rect 26236 38782 26350 38834
rect 26402 38782 26404 38834
rect 26236 38780 26404 38782
rect 26348 38770 26404 38780
rect 26460 38668 26516 41580
rect 26572 41412 26628 41422
rect 26572 40292 26628 41356
rect 26796 40516 26852 40526
rect 26684 40292 26740 40302
rect 26572 40290 26740 40292
rect 26572 40238 26686 40290
rect 26738 40238 26740 40290
rect 26572 40236 26740 40238
rect 26684 40226 26740 40236
rect 26796 39732 26852 40460
rect 25116 37998 25118 38050
rect 25170 37998 25172 38050
rect 25116 37986 25172 37998
rect 25228 38220 25620 38276
rect 25676 38388 25732 38398
rect 24780 37650 24836 37660
rect 25116 37604 25172 37614
rect 25116 37268 25172 37548
rect 25228 37492 25284 38220
rect 25340 38052 25396 38062
rect 25340 37958 25396 37996
rect 25564 37940 25620 37950
rect 25452 37938 25620 37940
rect 25452 37886 25566 37938
rect 25618 37886 25620 37938
rect 25452 37884 25620 37886
rect 25228 37436 25396 37492
rect 25228 37268 25284 37278
rect 25116 37266 25284 37268
rect 25116 37214 25230 37266
rect 25282 37214 25284 37266
rect 25116 37212 25284 37214
rect 25228 37202 25284 37212
rect 24332 36652 24612 36708
rect 25116 36708 25172 36718
rect 24108 34916 24164 35532
rect 24220 36036 24276 36046
rect 24220 35922 24276 35980
rect 24220 35870 24222 35922
rect 24274 35870 24276 35922
rect 24220 35026 24276 35870
rect 24220 34974 24222 35026
rect 24274 34974 24276 35026
rect 24220 34962 24276 34974
rect 23828 34188 23940 34244
rect 23996 34860 24164 34916
rect 23772 34178 23828 34188
rect 23436 33346 23492 33628
rect 23884 33906 23940 33918
rect 23884 33854 23886 33906
rect 23938 33854 23940 33906
rect 23884 33572 23940 33854
rect 23884 33506 23940 33516
rect 23436 33294 23438 33346
rect 23490 33294 23492 33346
rect 23436 33282 23492 33294
rect 23212 32946 23268 32956
rect 23324 33124 23380 33134
rect 23324 32562 23380 33068
rect 23660 33124 23716 33134
rect 23660 33030 23716 33068
rect 23884 32788 23940 32798
rect 23996 32788 24052 34860
rect 24332 34242 24388 36652
rect 25116 36614 25172 36652
rect 25340 36596 25396 37436
rect 25340 36530 25396 36540
rect 24444 36484 24500 36494
rect 24444 35924 24500 36428
rect 24556 36482 24612 36494
rect 24556 36430 24558 36482
rect 24610 36430 24612 36482
rect 24556 36372 24612 36430
rect 25452 36372 25508 37884
rect 25564 37874 25620 37884
rect 25564 37492 25620 37502
rect 25564 37378 25620 37436
rect 25564 37326 25566 37378
rect 25618 37326 25620 37378
rect 25564 37314 25620 37326
rect 24556 36306 24612 36316
rect 25004 36316 25508 36372
rect 25564 36932 25620 36942
rect 24444 35830 24500 35868
rect 24668 35698 24724 35710
rect 24668 35646 24670 35698
rect 24722 35646 24724 35698
rect 24556 35586 24612 35598
rect 24556 35534 24558 35586
rect 24610 35534 24612 35586
rect 24556 35028 24612 35534
rect 24668 35588 24724 35646
rect 24668 35522 24724 35532
rect 25004 35138 25060 36316
rect 25004 35086 25006 35138
rect 25058 35086 25060 35138
rect 25004 35074 25060 35086
rect 25116 36036 25172 36046
rect 24892 35028 24948 35038
rect 24556 35026 24948 35028
rect 24556 34974 24894 35026
rect 24946 34974 24948 35026
rect 24556 34972 24948 34974
rect 24892 34962 24948 34972
rect 24668 34580 24724 34590
rect 24332 34190 24334 34242
rect 24386 34190 24388 34242
rect 24332 34178 24388 34190
rect 24444 34244 24500 34254
rect 24444 34150 24500 34188
rect 24668 34242 24724 34524
rect 24668 34190 24670 34242
rect 24722 34190 24724 34242
rect 24668 34178 24724 34190
rect 24780 34132 24836 34142
rect 23884 32786 24052 32788
rect 23884 32734 23886 32786
rect 23938 32734 24052 32786
rect 23884 32732 24052 32734
rect 24108 33906 24164 33918
rect 24108 33854 24110 33906
rect 24162 33854 24164 33906
rect 24108 32788 24164 33854
rect 24668 33572 24724 33582
rect 24668 33458 24724 33516
rect 24668 33406 24670 33458
rect 24722 33406 24724 33458
rect 24668 33394 24724 33406
rect 24220 33348 24276 33358
rect 24220 33254 24276 33292
rect 23884 32722 23940 32732
rect 24108 32722 24164 32732
rect 24556 33234 24612 33246
rect 24556 33182 24558 33234
rect 24610 33182 24612 33234
rect 23324 32510 23326 32562
rect 23378 32510 23380 32562
rect 23324 32498 23380 32510
rect 24108 32564 24164 32574
rect 24556 32564 24612 33182
rect 24780 33122 24836 34076
rect 24780 33070 24782 33122
rect 24834 33070 24836 33122
rect 24668 32676 24724 32686
rect 24780 32676 24836 33070
rect 24724 32620 24836 32676
rect 24892 33796 24948 33806
rect 24668 32582 24724 32620
rect 24108 32562 24612 32564
rect 24108 32510 24110 32562
rect 24162 32510 24612 32562
rect 24108 32508 24612 32510
rect 24108 32452 24164 32508
rect 24108 32386 24164 32396
rect 24444 32002 24500 32014
rect 24444 31950 24446 32002
rect 24498 31950 24500 32002
rect 23996 31892 24052 31902
rect 24444 31892 24500 31950
rect 23772 31836 23996 31892
rect 23212 31668 23268 31678
rect 23660 31668 23716 31678
rect 23100 31666 23268 31668
rect 23100 31614 23214 31666
rect 23266 31614 23268 31666
rect 23100 31612 23268 31614
rect 23212 31602 23268 31612
rect 23548 31612 23660 31668
rect 22204 31166 22206 31218
rect 22258 31166 22260 31218
rect 22204 31154 22260 31166
rect 22876 31554 22932 31566
rect 22876 31502 22878 31554
rect 22930 31502 22932 31554
rect 21308 30942 21310 30994
rect 21362 30942 21364 30994
rect 21308 30930 21364 30942
rect 21756 30994 21812 31006
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 20972 30884 21028 30894
rect 19740 30772 19796 30782
rect 18732 30770 19796 30772
rect 18732 30718 19742 30770
rect 19794 30718 19796 30770
rect 18732 30716 19796 30718
rect 19740 30706 19796 30716
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18620 30146 18676 30158
rect 17724 30046 17726 30098
rect 17778 30046 17780 30098
rect 17052 28868 17108 28878
rect 16492 28866 17108 28868
rect 16492 28814 17054 28866
rect 17106 28814 17108 28866
rect 16492 28812 17108 28814
rect 17052 28802 17108 28812
rect 16380 28418 16436 28430
rect 16380 28366 16382 28418
rect 16434 28366 16436 28418
rect 16044 28084 16100 28094
rect 16044 27412 16100 28028
rect 15036 27188 15092 27198
rect 15036 26964 15092 27132
rect 14924 26962 15092 26964
rect 14924 26910 15038 26962
rect 15090 26910 15092 26962
rect 14924 26908 15092 26910
rect 14588 26852 14868 26908
rect 13468 26674 13524 26684
rect 14028 26516 14084 26526
rect 14028 26290 14084 26460
rect 14028 26238 14030 26290
rect 14082 26238 14084 26290
rect 14028 26226 14084 26238
rect 12348 25666 12404 25676
rect 14476 26068 14532 26078
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11340 25442 11396 25454
rect 14028 25506 14084 25518
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 12460 25284 12516 25294
rect 12460 25282 12628 25284
rect 12460 25230 12462 25282
rect 12514 25230 12628 25282
rect 12460 25228 12628 25230
rect 12460 25218 12516 25228
rect 12236 24612 12292 24622
rect 10444 24444 10836 24500
rect 9548 24050 9604 24062
rect 9548 23998 9550 24050
rect 9602 23998 9604 24050
rect 9100 23716 9156 23726
rect 8988 23660 9100 23716
rect 9100 23622 9156 23660
rect 9548 23380 9604 23998
rect 10444 24050 10500 24444
rect 10780 24388 10836 24444
rect 10780 24332 10948 24388
rect 10668 24276 10724 24286
rect 10724 24220 10836 24276
rect 10668 24210 10724 24220
rect 10444 23998 10446 24050
rect 10498 23998 10500 24050
rect 10444 23986 10500 23998
rect 9548 23314 9604 23324
rect 10108 23940 10164 23950
rect 8876 23202 8932 23212
rect 8988 23266 9044 23278
rect 8988 23214 8990 23266
rect 9042 23214 9044 23266
rect 8316 23062 8372 23100
rect 8540 23154 8820 23156
rect 8540 23102 8766 23154
rect 8818 23102 8820 23154
rect 8540 23100 8820 23102
rect 7980 22990 7982 23042
rect 8034 22990 8036 23042
rect 7980 21812 8036 22990
rect 8428 22148 8484 22158
rect 8428 22054 8484 22092
rect 8540 21924 8596 23100
rect 8764 23090 8820 23100
rect 7980 21746 8036 21756
rect 8316 21868 8596 21924
rect 8876 22482 8932 22494
rect 8876 22430 8878 22482
rect 8930 22430 8932 22482
rect 7980 20804 8036 20814
rect 7924 20802 8036 20804
rect 7924 20750 7982 20802
rect 8034 20750 8036 20802
rect 7924 20748 8036 20750
rect 7868 20710 7924 20748
rect 7980 20738 8036 20748
rect 7756 20578 7812 20590
rect 7756 20526 7758 20578
rect 7810 20526 7812 20578
rect 7756 20244 7812 20526
rect 8204 20244 8260 20254
rect 7756 20188 8148 20244
rect 8092 20130 8148 20188
rect 8092 20078 8094 20130
rect 8146 20078 8148 20130
rect 7980 20020 8036 20030
rect 7308 19966 7310 20018
rect 7362 19966 7364 20018
rect 7308 19954 7364 19966
rect 7532 20018 8036 20020
rect 7532 19966 7982 20018
rect 8034 19966 8036 20018
rect 7532 19964 8036 19966
rect 7532 19796 7588 19964
rect 7196 19740 7588 19796
rect 7644 19796 7700 19806
rect 7644 19702 7700 19740
rect 7420 19124 7476 19134
rect 7420 19030 7476 19068
rect 7868 18676 7924 18686
rect 7868 18582 7924 18620
rect 6972 18452 7028 18462
rect 6972 18358 7028 18396
rect 7196 18452 7252 18462
rect 7196 18358 7252 18396
rect 7420 18228 7476 18238
rect 7980 18228 8036 19964
rect 7308 18226 7476 18228
rect 7308 18174 7422 18226
rect 7474 18174 7476 18226
rect 7308 18172 7476 18174
rect 7308 17106 7364 18172
rect 7420 18162 7476 18172
rect 7868 18172 8036 18228
rect 7308 17054 7310 17106
rect 7362 17054 7364 17106
rect 6972 16884 7028 16894
rect 6972 16790 7028 16828
rect 7308 16772 7364 17054
rect 7084 16716 7308 16772
rect 7084 16098 7140 16716
rect 7308 16706 7364 16716
rect 7532 17668 7588 17678
rect 7084 16046 7086 16098
rect 7138 16046 7140 16098
rect 7084 16034 7140 16046
rect 6972 15988 7028 15998
rect 6972 15894 7028 15932
rect 7532 15988 7588 17612
rect 7644 16996 7700 17006
rect 7644 16902 7700 16940
rect 7756 16658 7812 16670
rect 7756 16606 7758 16658
rect 7810 16606 7812 16658
rect 7644 15988 7700 15998
rect 7532 15986 7700 15988
rect 7532 15934 7646 15986
rect 7698 15934 7700 15986
rect 7532 15932 7700 15934
rect 7084 15316 7140 15326
rect 7084 15148 7140 15260
rect 6860 15092 7028 15148
rect 7084 15092 7252 15148
rect 6748 14578 6804 14588
rect 6860 14868 6916 14878
rect 6636 14478 6638 14530
rect 6690 14478 6692 14530
rect 6412 14418 6468 14430
rect 6412 14366 6414 14418
rect 6466 14366 6468 14418
rect 6412 13636 6468 14366
rect 6524 13636 6580 13646
rect 6412 13580 6524 13636
rect 6524 13542 6580 13580
rect 6300 12964 6356 12974
rect 6300 12178 6356 12908
rect 6636 12964 6692 14478
rect 6748 13076 6804 13086
rect 6748 12982 6804 13020
rect 6636 12898 6692 12908
rect 6860 12292 6916 14812
rect 6972 14532 7028 15092
rect 6972 14476 7140 14532
rect 6972 14306 7028 14318
rect 6972 14254 6974 14306
rect 7026 14254 7028 14306
rect 6972 14084 7028 14254
rect 6972 14018 7028 14028
rect 7084 13860 7140 14476
rect 6300 12126 6302 12178
rect 6354 12126 6356 12178
rect 6300 12114 6356 12126
rect 6748 12236 6916 12292
rect 6972 13804 7140 13860
rect 6636 11170 6692 11182
rect 6636 11118 6638 11170
rect 6690 11118 6692 11170
rect 6636 10948 6692 11118
rect 6636 10882 6692 10892
rect 6076 10668 6468 10724
rect 5740 10558 5742 10610
rect 5794 10558 5796 10610
rect 5740 10546 5796 10558
rect 6188 10498 6244 10510
rect 6188 10446 6190 10498
rect 6242 10446 6244 10498
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 6076 10052 6132 10062
rect 5964 9940 6020 9950
rect 5964 9846 6020 9884
rect 3276 9538 3332 9548
rect 1708 9154 1764 9166
rect 1708 9102 1710 9154
rect 1762 9102 1764 9154
rect 1708 8820 1764 9102
rect 6076 9044 6132 9996
rect 6188 9268 6244 10446
rect 6412 9828 6468 10668
rect 6524 10612 6580 10622
rect 6524 10518 6580 10556
rect 6412 9772 6580 9828
rect 6188 9202 6244 9212
rect 6412 9602 6468 9614
rect 6412 9550 6414 9602
rect 6466 9550 6468 9602
rect 6188 9044 6244 9054
rect 6076 9042 6244 9044
rect 6076 8990 6190 9042
rect 6242 8990 6244 9042
rect 6076 8988 6244 8990
rect 6188 8978 6244 8988
rect 1708 8754 1764 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 6412 8484 6468 9550
rect 6412 8418 6468 8428
rect 6524 9266 6580 9772
rect 6524 9214 6526 9266
rect 6578 9214 6580 9266
rect 6300 8372 6356 8382
rect 6300 8278 6356 8316
rect 6524 8260 6580 9214
rect 6524 8194 6580 8204
rect 6748 8258 6804 12236
rect 6860 12068 6916 12078
rect 6860 11974 6916 12012
rect 6972 11396 7028 13804
rect 7196 13748 7252 15092
rect 7196 13682 7252 13692
rect 7308 14642 7364 14654
rect 7308 14590 7310 14642
rect 7362 14590 7364 14642
rect 7084 13634 7140 13646
rect 7084 13582 7086 13634
rect 7138 13582 7140 13634
rect 7084 13412 7140 13582
rect 7196 13524 7252 13534
rect 7196 13430 7252 13468
rect 7084 13346 7140 13356
rect 7084 12964 7140 12974
rect 7084 12870 7140 12908
rect 7308 12740 7364 14590
rect 7532 14642 7588 15932
rect 7644 15922 7700 15932
rect 7756 15428 7812 16606
rect 7644 14756 7700 14766
rect 7644 14662 7700 14700
rect 7532 14590 7534 14642
rect 7586 14590 7588 14642
rect 7532 14578 7588 14590
rect 7756 14532 7812 15372
rect 7868 16322 7924 18172
rect 7980 17668 8036 17678
rect 8092 17668 8148 20078
rect 8204 18676 8260 20188
rect 8204 18610 8260 18620
rect 8036 17612 8148 17668
rect 7980 17602 8036 17612
rect 7868 16270 7870 16322
rect 7922 16270 7924 16322
rect 7868 14868 7924 16270
rect 7980 17444 8036 17454
rect 7980 15092 8036 17388
rect 8316 16996 8372 21868
rect 8876 20580 8932 22430
rect 8988 22372 9044 23214
rect 8988 22306 9044 22316
rect 9324 23156 9380 23166
rect 9324 22370 9380 23100
rect 10108 23154 10164 23884
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 10108 23090 10164 23102
rect 10556 23156 10612 23166
rect 10556 23062 10612 23100
rect 9772 23044 9828 23054
rect 9772 23042 9940 23044
rect 9772 22990 9774 23042
rect 9826 22990 9940 23042
rect 9772 22988 9940 22990
rect 9772 22978 9828 22988
rect 9324 22318 9326 22370
rect 9378 22318 9380 22370
rect 9324 22306 9380 22318
rect 9660 22372 9716 22382
rect 9660 22278 9716 22316
rect 9772 22260 9828 22270
rect 9772 22166 9828 22204
rect 8876 20514 8932 20524
rect 9772 20580 9828 20590
rect 8652 20132 8708 20142
rect 8652 20038 8708 20076
rect 9660 19906 9716 19918
rect 9660 19854 9662 19906
rect 9714 19854 9716 19906
rect 8988 19234 9044 19246
rect 8988 19182 8990 19234
rect 9042 19182 9044 19234
rect 8652 19012 8708 19022
rect 8652 18674 8708 18956
rect 8652 18622 8654 18674
rect 8706 18622 8708 18674
rect 8652 18610 8708 18622
rect 8764 18452 8820 18462
rect 8428 17442 8484 17454
rect 8428 17390 8430 17442
rect 8482 17390 8484 17442
rect 8428 17108 8484 17390
rect 8484 17052 8708 17108
rect 8428 17014 8484 17052
rect 8316 16930 8372 16940
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 8428 16772 8484 16830
rect 8484 16716 8596 16772
rect 8428 16706 8484 16716
rect 8204 16324 8260 16334
rect 8204 16230 8260 16268
rect 8540 16098 8596 16716
rect 8540 16046 8542 16098
rect 8594 16046 8596 16098
rect 8540 16034 8596 16046
rect 8652 15876 8708 17052
rect 8428 15820 8708 15876
rect 8428 15204 8484 15820
rect 8428 15138 8484 15148
rect 8764 15314 8820 18396
rect 8876 17444 8932 17454
rect 8876 17350 8932 17388
rect 8988 17220 9044 19182
rect 9212 19122 9268 19134
rect 9212 19070 9214 19122
rect 9266 19070 9268 19122
rect 9212 19012 9268 19070
rect 9212 18946 9268 18956
rect 9660 19012 9716 19854
rect 9660 18946 9716 18956
rect 9772 19234 9828 20524
rect 9772 19182 9774 19234
rect 9826 19182 9828 19234
rect 9100 18900 9156 18910
rect 9100 18450 9156 18844
rect 9100 18398 9102 18450
rect 9154 18398 9156 18450
rect 9100 18386 9156 18398
rect 9548 18340 9604 18350
rect 9548 17666 9604 18284
rect 9660 18338 9716 18350
rect 9660 18286 9662 18338
rect 9714 18286 9716 18338
rect 9660 18116 9716 18286
rect 9660 18050 9716 18060
rect 9548 17614 9550 17666
rect 9602 17614 9604 17666
rect 9548 17602 9604 17614
rect 8764 15262 8766 15314
rect 8818 15262 8820 15314
rect 7980 15026 8036 15036
rect 8204 15092 8260 15102
rect 7868 14802 7924 14812
rect 7756 14530 8036 14532
rect 7756 14478 7758 14530
rect 7810 14478 8036 14530
rect 7756 14476 8036 14478
rect 7756 14466 7812 14476
rect 7980 13746 8036 14476
rect 8204 14084 8260 15036
rect 8316 15090 8372 15102
rect 8316 15038 8318 15090
rect 8370 15038 8372 15090
rect 8316 14980 8372 15038
rect 8316 14914 8372 14924
rect 8204 14018 8260 14028
rect 8316 14642 8372 14654
rect 8316 14590 8318 14642
rect 8370 14590 8372 14642
rect 7980 13694 7982 13746
rect 8034 13694 8036 13746
rect 7980 13682 8036 13694
rect 8092 13748 8148 13758
rect 7532 13634 7588 13646
rect 7532 13582 7534 13634
rect 7586 13582 7588 13634
rect 7532 13412 7588 13582
rect 7420 12852 7476 12862
rect 7420 12758 7476 12796
rect 6860 11340 7028 11396
rect 7084 12684 7364 12740
rect 6860 9828 6916 11340
rect 6972 11170 7028 11182
rect 6972 11118 6974 11170
rect 7026 11118 7028 11170
rect 6972 10948 7028 11118
rect 6972 10882 7028 10892
rect 7084 10836 7140 12684
rect 7532 12516 7588 13356
rect 7084 10742 7140 10780
rect 7196 12460 7588 12516
rect 7196 10500 7252 12460
rect 7308 12290 7364 12302
rect 7308 12238 7310 12290
rect 7362 12238 7364 12290
rect 7308 10948 7364 12238
rect 7532 12178 7588 12460
rect 7532 12126 7534 12178
rect 7586 12126 7588 12178
rect 7532 12114 7588 12126
rect 7644 13636 7700 13646
rect 7532 11508 7588 11518
rect 7532 11414 7588 11452
rect 7308 10882 7364 10892
rect 7532 10612 7588 10622
rect 7644 10612 7700 13580
rect 7868 12850 7924 12862
rect 7868 12798 7870 12850
rect 7922 12798 7924 12850
rect 7084 10444 7252 10500
rect 7420 10610 7700 10612
rect 7420 10558 7534 10610
rect 7586 10558 7700 10610
rect 7420 10556 7700 10558
rect 7756 10612 7812 10622
rect 6860 9772 7028 9828
rect 6860 9602 6916 9614
rect 6860 9550 6862 9602
rect 6914 9550 6916 9602
rect 6860 9492 6916 9550
rect 6860 9426 6916 9436
rect 6860 9268 6916 9278
rect 6860 9174 6916 9212
rect 6972 8596 7028 9772
rect 6748 8206 6750 8258
rect 6802 8206 6804 8258
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 6748 6916 6804 8206
rect 6748 6850 6804 6860
rect 6860 8540 7028 8596
rect 6860 7698 6916 8540
rect 6860 7646 6862 7698
rect 6914 7646 6916 7698
rect 6860 6914 6916 7646
rect 6860 6862 6862 6914
rect 6914 6862 6916 6914
rect 6860 6850 6916 6862
rect 7084 5908 7140 10444
rect 7420 10388 7476 10556
rect 7532 10546 7588 10556
rect 7196 10332 7476 10388
rect 7196 8258 7252 10332
rect 7756 9828 7812 10556
rect 7756 9734 7812 9772
rect 7868 9938 7924 12798
rect 8092 12740 8148 13692
rect 8204 13636 8260 13646
rect 8316 13636 8372 14590
rect 8540 14530 8596 14542
rect 8540 14478 8542 14530
rect 8594 14478 8596 14530
rect 8540 13972 8596 14478
rect 8540 13906 8596 13916
rect 8260 13580 8372 13636
rect 8428 13748 8484 13758
rect 8764 13748 8820 15262
rect 8428 13746 8820 13748
rect 8428 13694 8430 13746
rect 8482 13694 8820 13746
rect 8428 13692 8820 13694
rect 8876 17164 9044 17220
rect 9324 17442 9380 17454
rect 9324 17390 9326 17442
rect 9378 17390 9380 17442
rect 8204 13570 8260 13580
rect 8428 12852 8484 13692
rect 8428 12786 8484 12796
rect 8540 13524 8596 13534
rect 8540 12962 8596 13468
rect 8876 13412 8932 17164
rect 8988 16996 9044 17006
rect 8988 16902 9044 16940
rect 9324 16884 9380 17390
rect 9324 16818 9380 16828
rect 9772 16436 9828 19182
rect 9884 18452 9940 22988
rect 10780 22372 10836 24220
rect 10892 24052 10948 24332
rect 10892 24050 11172 24052
rect 10892 23998 10894 24050
rect 10946 23998 11172 24050
rect 10892 23996 11172 23998
rect 10892 23986 10948 23996
rect 11116 23156 11172 23996
rect 11900 24050 11956 24062
rect 11900 23998 11902 24050
rect 11954 23998 11956 24050
rect 11228 23940 11284 23950
rect 11228 23846 11284 23884
rect 11676 23492 11732 23502
rect 11564 23436 11676 23492
rect 11452 23156 11508 23166
rect 11116 23154 11508 23156
rect 11116 23102 11454 23154
rect 11506 23102 11508 23154
rect 11116 23100 11508 23102
rect 11004 23042 11060 23054
rect 11004 22990 11006 23042
rect 11058 22990 11060 23042
rect 10892 22484 10948 22494
rect 10892 22390 10948 22428
rect 10668 22316 10836 22372
rect 10220 22258 10276 22270
rect 10220 22206 10222 22258
rect 10274 22206 10276 22258
rect 10220 22148 10276 22206
rect 10220 22082 10276 22092
rect 10668 20804 10724 22316
rect 10780 22148 10836 22158
rect 10780 21810 10836 22092
rect 10780 21758 10782 21810
rect 10834 21758 10836 21810
rect 10780 21746 10836 21758
rect 10668 20748 10948 20804
rect 10668 20580 10724 20590
rect 10668 20486 10724 20524
rect 9996 20132 10052 20142
rect 9996 20018 10052 20076
rect 9996 19966 9998 20018
rect 10050 19966 10052 20018
rect 9996 19954 10052 19966
rect 10444 19908 10500 19918
rect 10556 19908 10612 19918
rect 10444 19906 10612 19908
rect 10444 19854 10446 19906
rect 10498 19854 10558 19906
rect 10610 19854 10612 19906
rect 10444 19852 10612 19854
rect 10108 19236 10164 19246
rect 10108 19142 10164 19180
rect 9884 18386 9940 18396
rect 10108 18338 10164 18350
rect 10108 18286 10110 18338
rect 10162 18286 10164 18338
rect 9996 17778 10052 17790
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9436 16380 9828 16436
rect 9884 17108 9940 17118
rect 9100 16098 9156 16110
rect 9100 16046 9102 16098
rect 9154 16046 9156 16098
rect 9100 14756 9156 16046
rect 9100 14690 9156 14700
rect 9212 14532 9268 14542
rect 9212 14438 9268 14476
rect 8876 13346 8932 13356
rect 8988 13634 9044 13646
rect 8988 13582 8990 13634
rect 9042 13582 9044 13634
rect 8540 12910 8542 12962
rect 8594 12910 8596 12962
rect 8092 12738 8260 12740
rect 8092 12686 8094 12738
rect 8146 12686 8260 12738
rect 8092 12684 8260 12686
rect 8092 12674 8148 12684
rect 7980 12180 8036 12190
rect 7980 12086 8036 12124
rect 7980 11170 8036 11182
rect 7980 11118 7982 11170
rect 8034 11118 8036 11170
rect 7980 10612 8036 11118
rect 8092 10948 8148 10958
rect 8092 10834 8148 10892
rect 8092 10782 8094 10834
rect 8146 10782 8148 10834
rect 8092 10770 8148 10782
rect 7980 10546 8036 10556
rect 7868 9886 7870 9938
rect 7922 9886 7924 9938
rect 7196 8206 7198 8258
rect 7250 8206 7252 8258
rect 7196 8194 7252 8206
rect 7308 9602 7364 9614
rect 7308 9550 7310 9602
rect 7362 9550 7364 9602
rect 7308 7924 7364 9550
rect 7868 9492 7924 9886
rect 7644 9436 7924 9492
rect 7420 8932 7476 8942
rect 7420 8930 7588 8932
rect 7420 8878 7422 8930
rect 7474 8878 7588 8930
rect 7420 8876 7588 8878
rect 7420 8866 7476 8876
rect 7308 7858 7364 7868
rect 7420 8484 7476 8494
rect 7196 7362 7252 7374
rect 7196 7310 7198 7362
rect 7250 7310 7252 7362
rect 7196 7250 7252 7310
rect 7196 7198 7198 7250
rect 7250 7198 7252 7250
rect 7196 7186 7252 7198
rect 7420 7250 7476 8428
rect 7420 7198 7422 7250
rect 7474 7198 7476 7250
rect 7420 7186 7476 7198
rect 7308 6914 7364 6926
rect 7308 6862 7310 6914
rect 7362 6862 7364 6914
rect 7308 6804 7364 6862
rect 7308 6710 7364 6748
rect 7196 5908 7252 5918
rect 7084 5852 7196 5908
rect 7196 5842 7252 5852
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 7532 5348 7588 8876
rect 7644 8372 7700 9436
rect 7756 9268 7812 9278
rect 7756 9042 7812 9212
rect 7868 9154 7924 9436
rect 7868 9102 7870 9154
rect 7922 9102 7924 9154
rect 7868 9090 7924 9102
rect 7756 8990 7758 9042
rect 7810 8990 7812 9042
rect 7756 8978 7812 8990
rect 8204 8820 8260 12684
rect 8428 12516 8484 12526
rect 8316 11956 8372 11966
rect 8316 11862 8372 11900
rect 8428 11506 8484 12460
rect 8428 11454 8430 11506
rect 8482 11454 8484 11506
rect 8428 11442 8484 11454
rect 8540 11060 8596 12910
rect 8988 11844 9044 13582
rect 9100 12404 9156 12414
rect 9100 12310 9156 12348
rect 8988 11778 9044 11788
rect 8428 11004 8596 11060
rect 8652 11506 8708 11518
rect 8652 11454 8654 11506
rect 8706 11454 8708 11506
rect 8428 9716 8484 11004
rect 8540 10836 8596 10846
rect 8540 10722 8596 10780
rect 8540 10670 8542 10722
rect 8594 10670 8596 10722
rect 8540 10658 8596 10670
rect 8652 10386 8708 11454
rect 8764 11508 8820 11518
rect 8764 11414 8820 11452
rect 9324 11172 9380 11182
rect 9324 11078 9380 11116
rect 8652 10334 8654 10386
rect 8706 10334 8708 10386
rect 8428 9660 8596 9716
rect 8316 9156 8372 9166
rect 8316 9062 8372 9100
rect 7644 8306 7700 8316
rect 7868 8764 8260 8820
rect 7644 8146 7700 8158
rect 7644 8094 7646 8146
rect 7698 8094 7700 8146
rect 7644 7252 7700 8094
rect 7644 6802 7700 7196
rect 7756 7362 7812 7374
rect 7756 7310 7758 7362
rect 7810 7310 7812 7362
rect 7756 7028 7812 7310
rect 7756 6962 7812 6972
rect 7644 6750 7646 6802
rect 7698 6750 7700 6802
rect 7644 6738 7700 6750
rect 7756 6244 7812 6254
rect 7756 6130 7812 6188
rect 7756 6078 7758 6130
rect 7810 6078 7812 6130
rect 7756 6066 7812 6078
rect 7532 5292 7812 5348
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 6972 3666 7028 3678
rect 6972 3614 6974 3666
rect 7026 3614 7028 3666
rect 6972 3388 7028 3614
rect 4844 3332 4900 3342
rect 5628 3332 5684 3342
rect 4732 3330 4900 3332
rect 4732 3278 4846 3330
rect 4898 3278 4900 3330
rect 4732 3276 4900 3278
rect 4732 800 4788 3276
rect 4844 3266 4900 3276
rect 5404 3330 5684 3332
rect 5404 3278 5630 3330
rect 5682 3278 5684 3330
rect 5404 3276 5684 3278
rect 5404 800 5460 3276
rect 5628 3266 5684 3276
rect 6748 3332 7028 3388
rect 7644 3332 7700 3342
rect 6748 800 6804 3332
rect 7420 3330 7700 3332
rect 7420 3278 7646 3330
rect 7698 3278 7700 3330
rect 7420 3276 7700 3278
rect 7420 800 7476 3276
rect 7644 3266 7700 3276
rect 7756 3332 7812 5292
rect 7756 3266 7812 3276
rect 7868 1428 7924 8764
rect 7980 8372 8036 8382
rect 7980 7698 8036 8316
rect 8428 8260 8484 8270
rect 7980 7646 7982 7698
rect 8034 7646 8036 7698
rect 7980 7634 8036 7646
rect 8092 8204 8428 8260
rect 7980 6804 8036 6814
rect 7980 6710 8036 6748
rect 8092 6130 8148 8204
rect 8428 8166 8484 8204
rect 8204 8036 8260 8046
rect 8540 8036 8596 9660
rect 8652 8708 8708 10334
rect 9436 10052 9492 16380
rect 9884 16324 9940 17052
rect 9660 16268 9940 16324
rect 9996 16322 10052 17726
rect 10108 16660 10164 18286
rect 10444 18116 10500 19852
rect 10556 19842 10612 19852
rect 10668 19796 10724 19806
rect 10668 19236 10724 19740
rect 10668 19234 10836 19236
rect 10668 19182 10670 19234
rect 10722 19182 10836 19234
rect 10668 19180 10836 19182
rect 10668 19170 10724 19180
rect 10780 18788 10836 19180
rect 10780 18722 10836 18732
rect 10556 18340 10612 18350
rect 10556 18246 10612 18284
rect 10444 18060 10612 18116
rect 10444 16884 10500 16894
rect 10108 16594 10164 16604
rect 10332 16658 10388 16670
rect 10332 16606 10334 16658
rect 10386 16606 10388 16658
rect 10332 16548 10388 16606
rect 10332 16482 10388 16492
rect 9996 16270 9998 16322
rect 10050 16270 10052 16322
rect 9548 15428 9604 15438
rect 9548 15334 9604 15372
rect 9548 14644 9604 14654
rect 9548 14530 9604 14588
rect 9548 14478 9550 14530
rect 9602 14478 9604 14530
rect 9548 14466 9604 14478
rect 9660 13972 9716 16268
rect 9884 16098 9940 16110
rect 9884 16046 9886 16098
rect 9938 16046 9940 16098
rect 9884 14532 9940 16046
rect 9996 15092 10052 16270
rect 10220 16324 10276 16334
rect 10444 16324 10500 16828
rect 10220 16322 10500 16324
rect 10220 16270 10222 16322
rect 10274 16270 10500 16322
rect 10220 16268 10500 16270
rect 10220 16258 10276 16268
rect 10444 15764 10500 15774
rect 10108 15428 10164 15438
rect 10108 15334 10164 15372
rect 10444 15426 10500 15708
rect 10444 15374 10446 15426
rect 10498 15374 10500 15426
rect 10444 15148 10500 15374
rect 9996 15026 10052 15036
rect 10332 15092 10500 15148
rect 10108 14756 10164 14766
rect 10164 14700 10276 14756
rect 10108 14690 10164 14700
rect 9884 14476 10164 14532
rect 9772 14420 9828 14430
rect 9772 14326 9828 14364
rect 9884 14308 9940 14318
rect 9884 14214 9940 14252
rect 9660 13916 9940 13972
rect 9772 13748 9828 13758
rect 9660 12852 9716 12862
rect 9660 12758 9716 12796
rect 9772 11618 9828 13692
rect 9884 12402 9940 13916
rect 10108 13076 10164 14476
rect 10220 14530 10276 14700
rect 10220 14478 10222 14530
rect 10274 14478 10276 14530
rect 10220 14466 10276 14478
rect 10332 14532 10388 15092
rect 10332 14466 10388 14476
rect 10444 14420 10500 14430
rect 10220 14196 10276 14206
rect 10220 13858 10276 14140
rect 10220 13806 10222 13858
rect 10274 13806 10276 13858
rect 10220 13794 10276 13806
rect 10444 13748 10500 14364
rect 10444 13682 10500 13692
rect 10108 13020 10276 13076
rect 10220 12964 10276 13020
rect 10220 12962 10500 12964
rect 10220 12910 10222 12962
rect 10274 12910 10500 12962
rect 10220 12908 10500 12910
rect 10220 12898 10276 12908
rect 10108 12852 10164 12862
rect 10108 12758 10164 12796
rect 9884 12350 9886 12402
rect 9938 12350 9940 12402
rect 9884 12338 9940 12350
rect 10332 12178 10388 12190
rect 10332 12126 10334 12178
rect 10386 12126 10388 12178
rect 10332 11844 10388 12126
rect 10332 11778 10388 11788
rect 9772 11566 9774 11618
rect 9826 11566 9828 11618
rect 9772 11554 9828 11566
rect 10108 11508 10164 11518
rect 10108 11414 10164 11452
rect 10332 11506 10388 11518
rect 10332 11454 10334 11506
rect 10386 11454 10388 11506
rect 10332 11396 10388 11454
rect 9436 9986 9492 9996
rect 9660 11170 9716 11182
rect 9660 11118 9662 11170
rect 9714 11118 9716 11170
rect 9660 11060 9716 11118
rect 8652 8642 8708 8652
rect 8876 9828 8932 9838
rect 8876 8258 8932 9772
rect 9436 9826 9492 9838
rect 9436 9774 9438 9826
rect 9490 9774 9492 9826
rect 9100 9492 9156 9502
rect 9100 9266 9156 9436
rect 9100 9214 9102 9266
rect 9154 9214 9156 9266
rect 9100 9202 9156 9214
rect 9436 9268 9492 9774
rect 9548 9268 9604 9278
rect 9492 9266 9604 9268
rect 9492 9214 9550 9266
rect 9602 9214 9604 9266
rect 9492 9212 9604 9214
rect 9436 9202 9492 9212
rect 9548 9202 9604 9212
rect 8876 8206 8878 8258
rect 8930 8206 8932 8258
rect 8876 8194 8932 8206
rect 9100 8372 9156 8382
rect 8204 8034 8372 8036
rect 8204 7982 8206 8034
rect 8258 7982 8372 8034
rect 8204 7980 8372 7982
rect 8204 7970 8260 7980
rect 8204 6916 8260 6926
rect 8204 6822 8260 6860
rect 8092 6078 8094 6130
rect 8146 6078 8148 6130
rect 8092 6066 8148 6078
rect 8316 2884 8372 7980
rect 8428 7980 8596 8036
rect 8428 6692 8484 7980
rect 9100 7698 9156 8316
rect 9548 8372 9604 8382
rect 9660 8372 9716 11004
rect 10108 10836 10164 10846
rect 10108 10742 10164 10780
rect 10332 10724 10388 11340
rect 10220 10722 10388 10724
rect 10220 10670 10334 10722
rect 10386 10670 10388 10722
rect 10220 10668 10388 10670
rect 9884 9940 9940 9950
rect 9884 9846 9940 9884
rect 9884 9716 9940 9726
rect 9884 9154 9940 9660
rect 9884 9102 9886 9154
rect 9938 9102 9940 9154
rect 9548 8370 9716 8372
rect 9548 8318 9550 8370
rect 9602 8318 9716 8370
rect 9548 8316 9716 8318
rect 9772 8596 9828 8606
rect 9548 8306 9604 8316
rect 9772 8260 9828 8540
rect 9884 8484 9940 9102
rect 10220 9154 10276 10668
rect 10332 10658 10388 10668
rect 10220 9102 10222 9154
rect 10274 9102 10276 9154
rect 10220 9090 10276 9102
rect 10444 9266 10500 12908
rect 10556 10052 10612 18060
rect 10668 17668 10724 17678
rect 10668 17574 10724 17612
rect 10780 16994 10836 17006
rect 10780 16942 10782 16994
rect 10834 16942 10836 16994
rect 10780 16324 10836 16942
rect 10668 15874 10724 15886
rect 10668 15822 10670 15874
rect 10722 15822 10724 15874
rect 10668 14980 10724 15822
rect 10780 15538 10836 16268
rect 10780 15486 10782 15538
rect 10834 15486 10836 15538
rect 10780 15474 10836 15486
rect 10892 15148 10948 20748
rect 11004 20692 11060 22990
rect 11228 22370 11284 22382
rect 11228 22318 11230 22370
rect 11282 22318 11284 22370
rect 11228 22148 11284 22318
rect 11228 22082 11284 22092
rect 11340 22370 11396 23100
rect 11452 23090 11508 23100
rect 11564 22596 11620 23436
rect 11676 23426 11732 23436
rect 11900 23380 11956 23998
rect 11340 22318 11342 22370
rect 11394 22318 11396 22370
rect 11116 21924 11172 21934
rect 11116 20914 11172 21868
rect 11116 20862 11118 20914
rect 11170 20862 11172 20914
rect 11116 20850 11172 20862
rect 11340 21476 11396 22318
rect 11004 20626 11060 20636
rect 11340 20018 11396 21420
rect 11340 19966 11342 20018
rect 11394 19966 11396 20018
rect 11004 19906 11060 19918
rect 11004 19854 11006 19906
rect 11058 19854 11060 19906
rect 11004 19796 11060 19854
rect 11004 19730 11060 19740
rect 11116 19796 11172 19806
rect 11340 19796 11396 19966
rect 11116 19794 11396 19796
rect 11116 19742 11118 19794
rect 11170 19742 11396 19794
rect 11116 19740 11396 19742
rect 11452 22540 11620 22596
rect 11676 22930 11732 22942
rect 11676 22878 11678 22930
rect 11730 22878 11732 22930
rect 11116 19730 11172 19740
rect 11116 19234 11172 19246
rect 11116 19182 11118 19234
rect 11170 19182 11172 19234
rect 11004 18676 11060 18686
rect 11116 18676 11172 19182
rect 11452 19012 11508 22540
rect 11564 22372 11620 22382
rect 11676 22372 11732 22878
rect 11620 22316 11732 22372
rect 11564 21586 11620 22316
rect 11788 22148 11844 22158
rect 11564 21534 11566 21586
rect 11618 21534 11620 21586
rect 11564 21522 11620 21534
rect 11676 22092 11788 22148
rect 11564 20692 11620 20702
rect 11564 20598 11620 20636
rect 11004 18674 11172 18676
rect 11004 18622 11006 18674
rect 11058 18622 11172 18674
rect 11004 18620 11172 18622
rect 11004 18610 11060 18620
rect 11116 18452 11172 18620
rect 11116 18386 11172 18396
rect 11228 18956 11508 19012
rect 11564 19012 11620 19022
rect 11116 17442 11172 17454
rect 11116 17390 11118 17442
rect 11170 17390 11172 17442
rect 11116 15876 11172 17390
rect 11228 15988 11284 18956
rect 11340 18788 11396 18798
rect 11340 17666 11396 18732
rect 11340 17614 11342 17666
rect 11394 17614 11396 17666
rect 11340 17602 11396 17614
rect 11452 18338 11508 18350
rect 11452 18286 11454 18338
rect 11506 18286 11508 18338
rect 11228 15922 11284 15932
rect 11116 15810 11172 15820
rect 11452 15148 11508 18286
rect 11564 16882 11620 18956
rect 11676 18452 11732 22092
rect 11788 22082 11844 22092
rect 11900 21924 11956 23324
rect 12012 23268 12068 23278
rect 12012 23174 12068 23212
rect 12124 22260 12180 22270
rect 12236 22260 12292 24556
rect 12572 23940 12628 25228
rect 12124 22258 12292 22260
rect 12124 22206 12126 22258
rect 12178 22206 12292 22258
rect 12124 22204 12292 22206
rect 12124 22194 12180 22204
rect 11900 21858 11956 21868
rect 12012 20578 12068 20590
rect 12012 20526 12014 20578
rect 12066 20526 12068 20578
rect 12012 20244 12068 20526
rect 12012 20178 12068 20188
rect 11900 19908 11956 19918
rect 11900 19814 11956 19852
rect 12124 19122 12180 19134
rect 12124 19070 12126 19122
rect 12178 19070 12180 19122
rect 12124 18564 12180 19070
rect 11900 18508 12180 18564
rect 11788 18452 11844 18462
rect 11732 18450 11844 18452
rect 11732 18398 11790 18450
rect 11842 18398 11844 18450
rect 11732 18396 11844 18398
rect 11676 18358 11732 18396
rect 11788 18386 11844 18396
rect 11900 18228 11956 18508
rect 12236 18228 12292 22204
rect 12348 23714 12404 23726
rect 12348 23662 12350 23714
rect 12402 23662 12404 23714
rect 12348 23380 12404 23662
rect 12460 23380 12516 23390
rect 12348 23378 12516 23380
rect 12348 23326 12462 23378
rect 12514 23326 12516 23378
rect 12348 23324 12516 23326
rect 12348 22148 12404 23324
rect 12460 23314 12516 23324
rect 12572 23266 12628 23884
rect 12572 23214 12574 23266
rect 12626 23214 12628 23266
rect 12572 23202 12628 23214
rect 12684 24610 12740 24622
rect 12684 24558 12686 24610
rect 12738 24558 12740 24610
rect 12684 23268 12740 24558
rect 13916 24612 13972 24622
rect 13916 24518 13972 24556
rect 13916 23940 13972 23950
rect 14028 23940 14084 25454
rect 14476 25506 14532 26012
rect 14476 25454 14478 25506
rect 14530 25454 14532 25506
rect 14476 25442 14532 25454
rect 14140 24724 14196 24734
rect 14140 24630 14196 24668
rect 13916 23938 14084 23940
rect 13916 23886 13918 23938
rect 13970 23886 14084 23938
rect 13916 23884 14084 23886
rect 14364 23940 14420 23950
rect 12796 23714 12852 23726
rect 12796 23662 12798 23714
rect 12850 23662 12852 23714
rect 12796 23380 12852 23662
rect 12796 23314 12852 23324
rect 13580 23380 13636 23390
rect 13580 23268 13636 23324
rect 13692 23268 13748 23278
rect 13580 23266 13748 23268
rect 13580 23214 13694 23266
rect 13746 23214 13748 23266
rect 13580 23212 13748 23214
rect 12684 23202 12740 23212
rect 13356 23156 13412 23166
rect 13020 23154 13412 23156
rect 13020 23102 13358 23154
rect 13410 23102 13412 23154
rect 13020 23100 13412 23102
rect 12908 23044 12964 23054
rect 12348 22082 12404 22092
rect 12572 22988 12908 23044
rect 12460 20916 12516 20926
rect 12460 20822 12516 20860
rect 12348 20132 12404 20142
rect 12348 20038 12404 20076
rect 11788 18172 11956 18228
rect 12124 18172 12292 18228
rect 12348 18676 12404 18686
rect 12348 18450 12404 18620
rect 12348 18398 12350 18450
rect 12402 18398 12404 18450
rect 12348 18340 12404 18398
rect 11564 16830 11566 16882
rect 11618 16830 11620 16882
rect 11564 16818 11620 16830
rect 11676 18116 11732 18126
rect 10892 15092 11172 15148
rect 10668 14924 10948 14980
rect 10668 14756 10724 14766
rect 10724 14700 10836 14756
rect 10668 14690 10724 14700
rect 10668 14418 10724 14430
rect 10668 14366 10670 14418
rect 10722 14366 10724 14418
rect 10668 14196 10724 14366
rect 10668 14130 10724 14140
rect 10668 13748 10724 13758
rect 10668 13654 10724 13692
rect 10668 11620 10724 11630
rect 10780 11620 10836 14700
rect 10892 12628 10948 14924
rect 11116 13636 11172 15092
rect 11228 15092 11508 15148
rect 11564 16212 11620 16222
rect 11676 16212 11732 18060
rect 11788 17108 11844 18172
rect 11900 17780 11956 17790
rect 11900 17686 11956 17724
rect 11900 17108 11956 17118
rect 11788 17052 11900 17108
rect 11900 17042 11956 17052
rect 12012 16996 12068 17006
rect 12012 16902 12068 16940
rect 11564 16210 11732 16212
rect 11564 16158 11566 16210
rect 11618 16158 11732 16210
rect 11564 16156 11732 16158
rect 12012 16212 12068 16222
rect 11228 14420 11284 15092
rect 11340 14868 11396 14878
rect 11340 14642 11396 14812
rect 11340 14590 11342 14642
rect 11394 14590 11396 14642
rect 11340 14578 11396 14590
rect 11228 14354 11284 14364
rect 11564 14196 11620 16156
rect 12012 16118 12068 16156
rect 11340 14140 11620 14196
rect 11676 15988 11732 15998
rect 11116 13634 11284 13636
rect 11116 13582 11118 13634
rect 11170 13582 11284 13634
rect 11116 13580 11284 13582
rect 11116 13570 11172 13580
rect 11116 12628 11172 12638
rect 10892 12572 11116 12628
rect 11116 12562 11172 12572
rect 10892 12292 10948 12302
rect 10892 12178 10948 12236
rect 10892 12126 10894 12178
rect 10946 12126 10948 12178
rect 10892 12114 10948 12126
rect 11004 12290 11060 12302
rect 11004 12238 11006 12290
rect 11058 12238 11060 12290
rect 11004 11788 11060 12238
rect 11116 12180 11172 12190
rect 11116 12066 11172 12124
rect 11116 12014 11118 12066
rect 11170 12014 11172 12066
rect 11116 12002 11172 12014
rect 10892 11732 11060 11788
rect 10892 11666 10948 11676
rect 10668 11618 10836 11620
rect 10668 11566 10670 11618
rect 10722 11566 10836 11618
rect 10668 11564 10836 11566
rect 10668 11554 10724 11564
rect 11116 11396 11172 11406
rect 10668 11284 10724 11322
rect 11116 11302 11172 11340
rect 10668 11218 10724 11228
rect 11228 11172 11284 13580
rect 11116 11116 11284 11172
rect 10556 9996 10724 10052
rect 10556 9828 10612 9838
rect 10556 9734 10612 9772
rect 10444 9214 10446 9266
rect 10498 9214 10500 9266
rect 10444 8708 10500 9214
rect 10556 8820 10612 8830
rect 10556 8726 10612 8764
rect 10108 8652 10500 8708
rect 9940 8428 10052 8484
rect 9884 8418 9940 8428
rect 9772 8194 9828 8204
rect 9884 8034 9940 8046
rect 9884 7982 9886 8034
rect 9938 7982 9940 8034
rect 9884 7924 9940 7982
rect 9884 7858 9940 7868
rect 9100 7646 9102 7698
rect 9154 7646 9156 7698
rect 9100 7634 9156 7646
rect 9548 7474 9604 7486
rect 9548 7422 9550 7474
rect 9602 7422 9604 7474
rect 8540 7364 8596 7374
rect 8540 7362 9044 7364
rect 8540 7310 8542 7362
rect 8594 7310 9044 7362
rect 8540 7308 9044 7310
rect 8540 7298 8596 7308
rect 8988 6916 9044 7308
rect 8988 6860 9492 6916
rect 9324 6692 9380 6702
rect 8428 6690 9380 6692
rect 8428 6638 9326 6690
rect 9378 6638 9380 6690
rect 8428 6636 9380 6638
rect 8428 6130 8484 6636
rect 9324 6626 9380 6636
rect 8428 6078 8430 6130
rect 8482 6078 8484 6130
rect 8428 6066 8484 6078
rect 8540 6466 8596 6478
rect 8540 6414 8542 6466
rect 8594 6414 8596 6466
rect 8540 5124 8596 6414
rect 8988 6468 9044 6478
rect 8988 6374 9044 6412
rect 9436 6020 9492 6860
rect 9548 6804 9604 7422
rect 9548 6738 9604 6748
rect 9884 6580 9940 6590
rect 9884 6486 9940 6524
rect 8540 5058 8596 5068
rect 8988 5794 9044 5806
rect 8988 5742 8990 5794
rect 9042 5742 9044 5794
rect 8988 3220 9044 5742
rect 9212 5236 9268 5246
rect 9212 5142 9268 5180
rect 9436 5012 9492 5964
rect 9660 6468 9716 6478
rect 9660 5234 9716 6412
rect 9772 6132 9828 6142
rect 9772 6038 9828 6076
rect 9660 5182 9662 5234
rect 9714 5182 9716 5234
rect 9660 5170 9716 5182
rect 9996 5012 10052 8428
rect 10108 7474 10164 8652
rect 10668 8260 10724 9996
rect 11004 9604 11060 9614
rect 11004 8930 11060 9548
rect 11004 8878 11006 8930
rect 11058 8878 11060 8930
rect 11004 8866 11060 8878
rect 10444 8204 10724 8260
rect 11004 8708 11060 8718
rect 10108 7422 10110 7474
rect 10162 7422 10164 7474
rect 10108 6692 10164 7422
rect 10332 8034 10388 8046
rect 10332 7982 10334 8034
rect 10386 7982 10388 8034
rect 10332 7252 10388 7982
rect 10332 7186 10388 7196
rect 10220 6692 10276 6702
rect 10108 6690 10276 6692
rect 10108 6638 10222 6690
rect 10274 6638 10276 6690
rect 10108 6636 10276 6638
rect 10220 6626 10276 6636
rect 10220 5908 10276 5918
rect 10108 5796 10164 5806
rect 10108 5234 10164 5740
rect 10108 5182 10110 5234
rect 10162 5182 10164 5234
rect 10108 5170 10164 5182
rect 10220 5124 10276 5852
rect 10332 5124 10388 5134
rect 10220 5122 10388 5124
rect 10220 5070 10334 5122
rect 10386 5070 10388 5122
rect 10220 5068 10388 5070
rect 10332 5058 10388 5068
rect 9436 4956 9828 5012
rect 9996 4956 10164 5012
rect 9772 4562 9828 4956
rect 9772 4510 9774 4562
rect 9826 4510 9828 4562
rect 9772 4498 9828 4510
rect 10108 4564 10164 4956
rect 10108 4498 10164 4508
rect 10444 4452 10500 8204
rect 10668 8034 10724 8046
rect 10668 7982 10670 8034
rect 10722 7982 10724 8034
rect 10668 7924 10724 7982
rect 11004 7924 11060 8652
rect 10668 7868 11060 7924
rect 10780 7364 10836 7374
rect 10780 7270 10836 7308
rect 10668 6692 10724 6702
rect 10668 6018 10724 6636
rect 10668 5966 10670 6018
rect 10722 5966 10724 6018
rect 10668 5954 10724 5966
rect 10780 6690 10836 6702
rect 10780 6638 10782 6690
rect 10834 6638 10836 6690
rect 10668 5572 10724 5582
rect 10668 5010 10724 5516
rect 10668 4958 10670 5010
rect 10722 4958 10724 5010
rect 10668 4946 10724 4958
rect 10332 4226 10388 4238
rect 10332 4174 10334 4226
rect 10386 4174 10388 4226
rect 10332 3778 10388 4174
rect 10332 3726 10334 3778
rect 10386 3726 10388 3778
rect 10332 3714 10388 3726
rect 10444 3666 10500 4396
rect 10444 3614 10446 3666
rect 10498 3614 10500 3666
rect 10444 3602 10500 3614
rect 10668 4564 10724 4574
rect 10668 3444 10724 4508
rect 10668 3378 10724 3388
rect 10780 3332 10836 6638
rect 10892 5124 10948 7868
rect 11116 7252 11172 11116
rect 11340 9828 11396 14140
rect 11564 13970 11620 13982
rect 11564 13918 11566 13970
rect 11618 13918 11620 13970
rect 11452 13748 11508 13758
rect 11452 13654 11508 13692
rect 11564 13188 11620 13918
rect 11452 12628 11508 12638
rect 11452 10724 11508 12572
rect 11564 12178 11620 13132
rect 11564 12126 11566 12178
rect 11618 12126 11620 12178
rect 11564 12068 11620 12126
rect 11564 12002 11620 12012
rect 11676 11844 11732 15932
rect 12124 15540 12180 18172
rect 12348 16996 12404 18284
rect 12348 16548 12404 16940
rect 12460 17666 12516 17678
rect 12460 17614 12462 17666
rect 12514 17614 12516 17666
rect 12460 16772 12516 17614
rect 12460 16706 12516 16716
rect 12348 16492 12516 16548
rect 12124 15484 12404 15540
rect 11788 15428 11844 15438
rect 11844 15372 12180 15428
rect 11788 15334 11844 15372
rect 11788 15092 11844 15102
rect 11788 14642 11844 15036
rect 11788 14590 11790 14642
rect 11842 14590 11844 14642
rect 11788 14578 11844 14590
rect 11900 14530 11956 14542
rect 11900 14478 11902 14530
rect 11954 14478 11956 14530
rect 11900 14196 11956 14478
rect 11900 14130 11956 14140
rect 12012 13858 12068 13870
rect 12012 13806 12014 13858
rect 12066 13806 12068 13858
rect 12012 13076 12068 13806
rect 11564 11788 11732 11844
rect 11900 13020 12012 13076
rect 11564 11394 11620 11788
rect 11564 11342 11566 11394
rect 11618 11342 11620 11394
rect 11564 10948 11620 11342
rect 11676 11284 11732 11294
rect 11676 11190 11732 11228
rect 11564 10882 11620 10892
rect 11676 10724 11732 10734
rect 11452 10668 11620 10724
rect 11340 9762 11396 9772
rect 11452 10052 11508 10062
rect 11228 9268 11284 9278
rect 11228 9042 11284 9212
rect 11228 8990 11230 9042
rect 11282 8990 11284 9042
rect 11228 8978 11284 8990
rect 11452 8930 11508 9996
rect 11452 8878 11454 8930
rect 11506 8878 11508 8930
rect 11228 8260 11284 8270
rect 11228 8166 11284 8204
rect 11340 7700 11396 7710
rect 11340 7362 11396 7644
rect 11340 7310 11342 7362
rect 11394 7310 11396 7362
rect 11116 7196 11284 7252
rect 11116 6692 11172 6702
rect 11116 6598 11172 6636
rect 11228 6130 11284 7196
rect 11340 6356 11396 7310
rect 11340 6290 11396 6300
rect 11452 7140 11508 8878
rect 11452 6804 11508 7084
rect 11564 7028 11620 10668
rect 11676 9714 11732 10668
rect 11676 9662 11678 9714
rect 11730 9662 11732 9714
rect 11676 7476 11732 9662
rect 11788 10500 11844 10510
rect 11788 7924 11844 10444
rect 11900 9044 11956 13020
rect 12012 13010 12068 13020
rect 12124 12962 12180 15372
rect 12348 15148 12404 15484
rect 12460 15314 12516 16492
rect 12572 16210 12628 22988
rect 12908 22978 12964 22988
rect 13020 22484 13076 23100
rect 13356 23090 13412 23100
rect 12908 22148 12964 22158
rect 12908 22054 12964 22092
rect 12684 21474 12740 21486
rect 12684 21422 12686 21474
rect 12738 21422 12740 21474
rect 12684 20020 12740 21422
rect 12908 20804 12964 20814
rect 13020 20804 13076 22428
rect 13468 22148 13524 22158
rect 13244 21476 13300 21486
rect 13244 21382 13300 21420
rect 13468 20916 13524 22092
rect 12908 20802 13076 20804
rect 12908 20750 12910 20802
rect 12962 20750 13076 20802
rect 12908 20748 13076 20750
rect 13244 20860 13468 20916
rect 12908 20738 12964 20748
rect 13132 20020 13188 20030
rect 12684 20018 13188 20020
rect 12684 19966 13134 20018
rect 13186 19966 13188 20018
rect 12684 19964 13188 19966
rect 12908 19012 12964 19050
rect 12908 18946 12964 18956
rect 12908 18788 12964 18798
rect 12796 18564 12852 18574
rect 12796 18450 12852 18508
rect 12796 18398 12798 18450
rect 12850 18398 12852 18450
rect 12796 18386 12852 18398
rect 12908 17778 12964 18732
rect 13132 18564 13188 19964
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17714 12964 17726
rect 13020 18562 13188 18564
rect 13020 18510 13134 18562
rect 13186 18510 13188 18562
rect 13020 18508 13188 18510
rect 13020 17556 13076 18508
rect 13132 18498 13188 18508
rect 12572 16158 12574 16210
rect 12626 16158 12628 16210
rect 12572 16146 12628 16158
rect 12908 16436 12964 16446
rect 12908 16210 12964 16380
rect 12908 16158 12910 16210
rect 12962 16158 12964 16210
rect 12908 16146 12964 16158
rect 12460 15262 12462 15314
rect 12514 15262 12516 15314
rect 12460 15250 12516 15262
rect 12684 15426 12740 15438
rect 12684 15374 12686 15426
rect 12738 15374 12740 15426
rect 12124 12910 12126 12962
rect 12178 12910 12180 12962
rect 12124 12292 12180 12910
rect 12236 15092 12404 15148
rect 12236 12628 12292 15092
rect 12684 14196 12740 15374
rect 12796 15314 12852 15326
rect 12796 15262 12798 15314
rect 12850 15262 12852 15314
rect 12796 15092 12852 15262
rect 12796 15026 12852 15036
rect 12684 14130 12740 14140
rect 12796 14642 12852 14654
rect 12796 14590 12798 14642
rect 12850 14590 12852 14642
rect 12796 13860 12852 14590
rect 13020 14530 13076 17500
rect 13244 15148 13300 20860
rect 13468 20850 13524 20860
rect 13580 20578 13636 20590
rect 13580 20526 13582 20578
rect 13634 20526 13636 20578
rect 13580 20468 13636 20526
rect 13580 20402 13636 20412
rect 13692 20244 13748 23212
rect 13916 23156 13972 23884
rect 13804 22372 13860 22382
rect 13916 22372 13972 23100
rect 13804 22370 13916 22372
rect 13804 22318 13806 22370
rect 13858 22318 13916 22370
rect 13804 22316 13916 22318
rect 13804 22306 13860 22316
rect 13916 22278 13972 22316
rect 14252 22370 14308 22382
rect 14252 22318 14254 22370
rect 14306 22318 14308 22370
rect 14252 21812 14308 22318
rect 14252 21746 14308 21756
rect 14140 21586 14196 21598
rect 14140 21534 14142 21586
rect 14194 21534 14196 21586
rect 13804 21474 13860 21486
rect 13804 21422 13806 21474
rect 13858 21422 13860 21474
rect 13804 20916 13860 21422
rect 13804 20850 13860 20860
rect 14028 20804 14084 20814
rect 14140 20804 14196 21534
rect 14028 20802 14196 20804
rect 14028 20750 14030 20802
rect 14082 20750 14196 20802
rect 14028 20748 14196 20750
rect 14028 20356 14084 20748
rect 14028 20290 14084 20300
rect 13692 20188 13972 20244
rect 13692 19234 13748 19246
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13580 19122 13636 19134
rect 13580 19070 13582 19122
rect 13634 19070 13636 19122
rect 13580 17780 13636 19070
rect 13692 18676 13748 19182
rect 13692 18610 13748 18620
rect 13692 18452 13748 18462
rect 13692 18358 13748 18396
rect 13580 17668 13636 17724
rect 13804 18338 13860 18350
rect 13804 18286 13806 18338
rect 13858 18286 13860 18338
rect 13580 17612 13748 17668
rect 13580 17442 13636 17454
rect 13580 17390 13582 17442
rect 13634 17390 13636 17442
rect 13356 16882 13412 16894
rect 13356 16830 13358 16882
rect 13410 16830 13412 16882
rect 13356 16772 13412 16830
rect 13468 16772 13524 16782
rect 13356 16716 13468 16772
rect 13468 16706 13524 16716
rect 13468 16548 13524 16558
rect 13020 14478 13022 14530
rect 13074 14478 13076 14530
rect 13020 14466 13076 14478
rect 13132 15092 13300 15148
rect 13356 16212 13412 16222
rect 12796 13794 12852 13804
rect 13020 13972 13076 13982
rect 12908 13076 12964 13086
rect 13020 13076 13076 13916
rect 12908 13074 13076 13076
rect 12908 13022 12910 13074
rect 12962 13022 13076 13074
rect 12908 13020 13076 13022
rect 12908 13010 12964 13020
rect 12348 12740 12404 12750
rect 12348 12646 12404 12684
rect 12236 12404 12292 12572
rect 12236 12338 12292 12348
rect 12572 12404 12628 12414
rect 12012 12068 12068 12078
rect 12012 11844 12068 12012
rect 12012 10610 12068 11788
rect 12124 11394 12180 12236
rect 12124 11342 12126 11394
rect 12178 11342 12180 11394
rect 12124 11330 12180 11342
rect 12460 12290 12516 12302
rect 12460 12238 12462 12290
rect 12514 12238 12516 12290
rect 12012 10558 12014 10610
rect 12066 10558 12068 10610
rect 12012 10546 12068 10558
rect 12124 10612 12180 10622
rect 11900 8370 11956 8988
rect 11900 8318 11902 8370
rect 11954 8318 11956 8370
rect 11900 8306 11956 8318
rect 11788 7858 11844 7868
rect 11788 7476 11844 7486
rect 11676 7474 11844 7476
rect 11676 7422 11790 7474
rect 11842 7422 11844 7474
rect 11676 7420 11844 7422
rect 11676 7028 11732 7038
rect 11564 6972 11676 7028
rect 11676 6962 11732 6972
rect 11228 6078 11230 6130
rect 11282 6078 11284 6130
rect 11228 6066 11284 6078
rect 11116 5124 11172 5134
rect 10892 5122 11172 5124
rect 10892 5070 11118 5122
rect 11170 5070 11172 5122
rect 10892 5068 11172 5070
rect 11116 5058 11172 5068
rect 10892 4564 10948 4574
rect 10892 3666 10948 4508
rect 11228 4564 11284 4574
rect 11452 4564 11508 6748
rect 11676 6804 11732 6814
rect 11676 6130 11732 6748
rect 11788 6690 11844 7420
rect 11788 6638 11790 6690
rect 11842 6638 11844 6690
rect 11788 6626 11844 6638
rect 11676 6078 11678 6130
rect 11730 6078 11732 6130
rect 11676 6066 11732 6078
rect 12124 6132 12180 10556
rect 12348 10610 12404 10622
rect 12348 10558 12350 10610
rect 12402 10558 12404 10610
rect 12236 9828 12292 9838
rect 12236 9734 12292 9772
rect 12348 9604 12404 10558
rect 12460 10164 12516 12238
rect 12572 12066 12628 12348
rect 12684 12180 12740 12190
rect 12684 12086 12740 12124
rect 12572 12014 12574 12066
rect 12626 12014 12628 12066
rect 12572 12002 12628 12014
rect 12572 11732 12628 11742
rect 12572 11506 12628 11676
rect 12572 11454 12574 11506
rect 12626 11454 12628 11506
rect 12572 11396 12628 11454
rect 12572 11330 12628 11340
rect 12908 10724 12964 10734
rect 12908 10630 12964 10668
rect 12460 10098 12516 10108
rect 12908 9828 12964 9838
rect 12908 9734 12964 9772
rect 12684 9716 12740 9726
rect 12684 9622 12740 9660
rect 12404 9548 12628 9604
rect 12348 9538 12404 9548
rect 12572 9268 12628 9548
rect 12796 9602 12852 9614
rect 12796 9550 12798 9602
rect 12850 9550 12852 9602
rect 12572 9212 12740 9268
rect 12572 9044 12628 9054
rect 12572 8950 12628 8988
rect 12348 8708 12404 8718
rect 12236 8260 12292 8270
rect 12236 8166 12292 8204
rect 12124 5908 12180 6076
rect 12236 6132 12292 6142
rect 12348 6132 12404 8652
rect 12684 7586 12740 9212
rect 12796 9156 12852 9550
rect 12796 9090 12852 9100
rect 12908 8484 12964 8494
rect 13020 8484 13076 13020
rect 13132 10164 13188 15092
rect 13244 14196 13300 14206
rect 13244 13746 13300 14140
rect 13244 13694 13246 13746
rect 13298 13694 13300 13746
rect 13244 13682 13300 13694
rect 13244 12180 13300 12190
rect 13356 12180 13412 16156
rect 13468 16098 13524 16492
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 16034 13524 16046
rect 13580 15148 13636 17390
rect 13692 15652 13748 17612
rect 13804 16996 13860 18286
rect 13916 17666 13972 20188
rect 14364 19796 14420 23884
rect 14588 23940 14644 23950
rect 14588 23042 14644 23884
rect 14812 23380 14868 26852
rect 14924 26628 14980 26908
rect 15036 26898 15092 26908
rect 16044 26962 16100 27356
rect 16044 26910 16046 26962
rect 16098 26910 16100 26962
rect 16044 26898 16100 26910
rect 16268 26964 16324 26974
rect 15260 26852 15316 26862
rect 15260 26850 15540 26852
rect 15260 26798 15262 26850
rect 15314 26798 15540 26850
rect 15260 26796 15540 26798
rect 15260 26786 15316 26796
rect 14924 26562 14980 26572
rect 15036 26068 15092 26078
rect 15092 26012 15316 26068
rect 15036 25974 15092 26012
rect 15260 25618 15316 26012
rect 15260 25566 15262 25618
rect 15314 25566 15316 25618
rect 15260 25554 15316 25566
rect 15372 25396 15428 25406
rect 14924 24724 14980 24734
rect 14924 23938 14980 24668
rect 15260 24722 15316 24734
rect 15260 24670 15262 24722
rect 15314 24670 15316 24722
rect 15260 24612 15316 24670
rect 15260 24546 15316 24556
rect 14924 23886 14926 23938
rect 14978 23886 14980 23938
rect 14924 23874 14980 23886
rect 15372 23938 15428 25340
rect 15484 24948 15540 26796
rect 16268 25732 16324 26908
rect 16380 26516 16436 28366
rect 17724 27972 17780 30046
rect 18284 30100 18340 30110
rect 18284 30006 18340 30044
rect 18732 30100 18788 30110
rect 18732 30006 18788 30044
rect 18956 30100 19012 30110
rect 18956 30006 19012 30044
rect 19180 30098 19236 30110
rect 19180 30046 19182 30098
rect 19234 30046 19236 30098
rect 19068 29988 19124 29998
rect 18956 29314 19012 29326
rect 18956 29262 18958 29314
rect 19010 29262 19012 29314
rect 18396 29204 18452 29214
rect 18396 28530 18452 29148
rect 18956 29092 19012 29262
rect 18396 28478 18398 28530
rect 18450 28478 18452 28530
rect 18396 28466 18452 28478
rect 18508 28532 18564 28542
rect 18508 28438 18564 28476
rect 18732 28418 18788 28430
rect 18732 28366 18734 28418
rect 18786 28366 18788 28418
rect 17948 27972 18004 27982
rect 17724 27916 17948 27972
rect 17948 27878 18004 27916
rect 18620 27972 18676 27982
rect 18732 27972 18788 28366
rect 18620 27970 18788 27972
rect 18620 27918 18622 27970
rect 18674 27918 18788 27970
rect 18620 27916 18788 27918
rect 18620 27906 18676 27916
rect 16380 26450 16436 26460
rect 18172 27858 18228 27870
rect 18172 27806 18174 27858
rect 18226 27806 18228 27858
rect 16268 25666 16324 25676
rect 17836 25508 17892 25518
rect 17836 25414 17892 25452
rect 18172 25508 18228 27806
rect 18844 27860 18900 27870
rect 18844 27766 18900 27804
rect 18732 27636 18788 27646
rect 18732 27542 18788 27580
rect 18732 27188 18788 27198
rect 18956 27188 19012 29036
rect 19068 29202 19124 29932
rect 19068 29150 19070 29202
rect 19122 29150 19124 29202
rect 19068 28980 19124 29150
rect 19180 29204 19236 30046
rect 19628 30100 19684 30110
rect 19628 30006 19684 30044
rect 20412 30100 20468 30110
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19180 29138 19236 29148
rect 19628 29650 19684 29662
rect 19628 29598 19630 29650
rect 19682 29598 19684 29650
rect 19068 28914 19124 28924
rect 18788 27132 19012 27188
rect 19068 28532 19124 28542
rect 19068 28420 19124 28476
rect 19180 28420 19236 28430
rect 19068 28418 19236 28420
rect 19068 28366 19182 28418
rect 19234 28366 19236 28418
rect 19068 28364 19236 28366
rect 18396 27076 18452 27086
rect 18396 26982 18452 27020
rect 18732 27074 18788 27132
rect 18732 27022 18734 27074
rect 18786 27022 18788 27074
rect 18732 27010 18788 27022
rect 19068 26908 19124 28364
rect 19180 28354 19236 28364
rect 19628 28084 19684 29598
rect 20412 28642 20468 30044
rect 20972 29988 21028 30828
rect 21756 30884 21812 30942
rect 21756 30324 21812 30828
rect 22316 30884 22372 30894
rect 22316 30790 22372 30828
rect 22764 30884 22820 30894
rect 22876 30884 22932 31502
rect 23436 31220 23492 31230
rect 23436 31126 23492 31164
rect 23548 31218 23604 31612
rect 23660 31602 23716 31612
rect 23548 31166 23550 31218
rect 23602 31166 23604 31218
rect 23548 31154 23604 31166
rect 23772 31218 23828 31836
rect 23996 31798 24052 31836
rect 24108 31836 24500 31892
rect 23772 31166 23774 31218
rect 23826 31166 23828 31218
rect 23772 31154 23828 31166
rect 23884 31108 23940 31118
rect 24108 31108 24164 31836
rect 23884 31106 24164 31108
rect 23884 31054 23886 31106
rect 23938 31054 24164 31106
rect 23884 31052 24164 31054
rect 24332 31666 24388 31678
rect 24332 31614 24334 31666
rect 24386 31614 24388 31666
rect 23884 31042 23940 31052
rect 24220 30996 24276 31006
rect 24332 30996 24388 31614
rect 24444 31554 24500 31566
rect 24444 31502 24446 31554
rect 24498 31502 24500 31554
rect 24444 31444 24500 31502
rect 24780 31444 24836 31454
rect 24444 31388 24780 31444
rect 24444 31220 24500 31230
rect 24444 31126 24500 31164
rect 24668 31218 24724 31388
rect 24780 31378 24836 31388
rect 24668 31166 24670 31218
rect 24722 31166 24724 31218
rect 24668 31154 24724 31166
rect 24892 31220 24948 33740
rect 25116 31668 25172 35980
rect 25340 35700 25396 35710
rect 25340 35606 25396 35644
rect 25564 35698 25620 36876
rect 25564 35646 25566 35698
rect 25618 35646 25620 35698
rect 25564 35364 25620 35646
rect 25564 35298 25620 35308
rect 25452 34692 25508 34702
rect 25452 34132 25508 34636
rect 25452 34066 25508 34076
rect 25564 34018 25620 34030
rect 25564 33966 25566 34018
rect 25618 33966 25620 34018
rect 25564 33908 25620 33966
rect 25228 33852 25620 33908
rect 25228 32900 25284 33852
rect 25676 33796 25732 38332
rect 26012 38162 26068 38174
rect 26012 38110 26014 38162
rect 26066 38110 26068 38162
rect 26012 38052 26068 38110
rect 26012 37986 26068 37996
rect 26124 38050 26180 38668
rect 26124 37998 26126 38050
rect 26178 37998 26180 38050
rect 26124 37986 26180 37998
rect 26236 38612 26516 38668
rect 26572 39676 26852 39732
rect 26908 40292 26964 43036
rect 27020 42868 27076 42878
rect 27020 42866 27188 42868
rect 27020 42814 27022 42866
rect 27074 42814 27188 42866
rect 27020 42812 27188 42814
rect 27020 42802 27076 42812
rect 27020 42644 27076 42654
rect 27020 41972 27076 42588
rect 27132 42420 27188 42812
rect 27132 42354 27188 42364
rect 27356 42196 27412 43036
rect 27468 42868 27524 42878
rect 27468 42532 27524 42812
rect 27916 42644 27972 45388
rect 28028 45330 28084 45388
rect 28028 45278 28030 45330
rect 28082 45278 28084 45330
rect 28028 45266 28084 45278
rect 28140 45108 28196 45612
rect 28028 45052 28196 45108
rect 28028 44996 28084 45052
rect 28028 43652 28084 44940
rect 28140 44884 28196 44894
rect 28140 44790 28196 44828
rect 28252 44324 28308 44334
rect 28252 44230 28308 44268
rect 28028 43596 28308 43652
rect 28140 43426 28196 43438
rect 28140 43374 28142 43426
rect 28194 43374 28196 43426
rect 28140 43316 28196 43374
rect 28140 43250 28196 43260
rect 28140 42868 28196 42878
rect 28140 42774 28196 42812
rect 27468 42466 27524 42476
rect 27580 42588 27972 42644
rect 28140 42644 28196 42654
rect 27356 42082 27412 42140
rect 27356 42030 27358 42082
rect 27410 42030 27412 42082
rect 27356 42018 27412 42030
rect 27468 42308 27524 42318
rect 27020 41970 27300 41972
rect 27020 41918 27022 41970
rect 27074 41918 27300 41970
rect 27020 41916 27300 41918
rect 27020 41906 27076 41916
rect 27020 41300 27076 41310
rect 27020 41186 27076 41244
rect 27020 41134 27022 41186
rect 27074 41134 27076 41186
rect 27020 41122 27076 41134
rect 27244 40626 27300 41916
rect 27468 41524 27524 42252
rect 27244 40574 27246 40626
rect 27298 40574 27300 40626
rect 27244 40562 27300 40574
rect 27356 41468 27524 41524
rect 27356 40404 27412 41468
rect 27468 41300 27524 41310
rect 27580 41300 27636 42588
rect 27916 42194 27972 42206
rect 27916 42142 27918 42194
rect 27970 42142 27972 42194
rect 27916 41972 27972 42142
rect 27916 41906 27972 41916
rect 28028 41970 28084 41982
rect 28028 41918 28030 41970
rect 28082 41918 28084 41970
rect 28028 41748 28084 41918
rect 28028 41682 28084 41692
rect 28140 41412 28196 42588
rect 28140 41346 28196 41356
rect 27468 41298 27580 41300
rect 27468 41246 27470 41298
rect 27522 41246 27580 41298
rect 27468 41244 27580 41246
rect 27468 41234 27524 41244
rect 27580 41206 27636 41244
rect 28028 41188 28084 41198
rect 28028 41094 28084 41132
rect 27468 40628 27524 40638
rect 27468 40626 27860 40628
rect 27468 40574 27470 40626
rect 27522 40574 27860 40626
rect 27468 40572 27860 40574
rect 27468 40562 27524 40572
rect 27580 40404 27636 40414
rect 27356 40402 27636 40404
rect 27356 40350 27582 40402
rect 27634 40350 27636 40402
rect 27356 40348 27636 40350
rect 27580 40338 27636 40348
rect 27020 40292 27076 40302
rect 26908 40290 27076 40292
rect 26908 40238 27022 40290
rect 27074 40238 27076 40290
rect 26908 40236 27076 40238
rect 26572 38836 26628 39676
rect 26908 39620 26964 40236
rect 27020 40226 27076 40236
rect 25900 37940 25956 37950
rect 25900 37846 25956 37884
rect 26012 36484 26068 36494
rect 26012 36390 26068 36428
rect 26236 35586 26292 38612
rect 26348 37826 26404 37838
rect 26348 37774 26350 37826
rect 26402 37774 26404 37826
rect 26348 37716 26404 37774
rect 26348 37154 26404 37660
rect 26348 37102 26350 37154
rect 26402 37102 26404 37154
rect 26348 37090 26404 37102
rect 26572 36596 26628 38780
rect 26684 39564 26964 39620
rect 27356 39956 27412 39966
rect 27356 39618 27412 39900
rect 27580 39620 27636 39630
rect 27356 39566 27358 39618
rect 27410 39566 27412 39618
rect 26684 38948 26740 39564
rect 27356 39554 27412 39566
rect 27468 39618 27636 39620
rect 27468 39566 27582 39618
rect 27634 39566 27636 39618
rect 27468 39564 27636 39566
rect 26908 39394 26964 39406
rect 26908 39342 26910 39394
rect 26962 39342 26964 39394
rect 26908 39284 26964 39342
rect 27468 39284 27524 39564
rect 27580 39554 27636 39564
rect 26908 39228 27524 39284
rect 26684 37716 26740 38892
rect 26908 38500 26964 38510
rect 26684 37650 26740 37660
rect 26796 37826 26852 37838
rect 26796 37774 26798 37826
rect 26850 37774 26852 37826
rect 26796 37380 26852 37774
rect 26796 37314 26852 37324
rect 26908 37268 26964 38444
rect 26908 37156 26964 37212
rect 26572 36530 26628 36540
rect 26796 37100 26964 37156
rect 27020 37266 27076 37278
rect 27020 37214 27022 37266
rect 27074 37214 27076 37266
rect 26796 36594 26852 37100
rect 27020 37044 27076 37214
rect 26796 36542 26798 36594
rect 26850 36542 26852 36594
rect 26796 36530 26852 36542
rect 26908 36988 27076 37044
rect 26796 36260 26852 36270
rect 26236 35534 26238 35586
rect 26290 35534 26292 35586
rect 26236 35522 26292 35534
rect 26572 35924 26628 35934
rect 26236 35252 26292 35262
rect 25788 34916 25844 34926
rect 25788 34822 25844 34860
rect 26012 34914 26068 34926
rect 26012 34862 26014 34914
rect 26066 34862 26068 34914
rect 25900 34580 25956 34590
rect 25676 33730 25732 33740
rect 25788 34468 25844 34478
rect 25676 33572 25732 33582
rect 25676 33478 25732 33516
rect 25340 33460 25396 33470
rect 25340 33366 25396 33404
rect 25228 32834 25284 32844
rect 25452 33346 25508 33358
rect 25452 33294 25454 33346
rect 25506 33294 25508 33346
rect 25452 32788 25508 33294
rect 25788 32900 25844 34412
rect 25452 32722 25508 32732
rect 25564 32844 25844 32900
rect 25452 32564 25508 32574
rect 25564 32564 25620 32844
rect 25900 32786 25956 34524
rect 26012 34244 26068 34862
rect 26012 34178 26068 34188
rect 26124 34130 26180 34142
rect 26124 34078 26126 34130
rect 26178 34078 26180 34130
rect 26124 34020 26180 34078
rect 26124 33954 26180 33964
rect 26236 33458 26292 35196
rect 26348 34690 26404 34702
rect 26348 34638 26350 34690
rect 26402 34638 26404 34690
rect 26348 34132 26404 34638
rect 26348 34066 26404 34076
rect 26236 33406 26238 33458
rect 26290 33406 26292 33458
rect 26236 33394 26292 33406
rect 26572 34018 26628 35868
rect 26684 35698 26740 35710
rect 26684 35646 26686 35698
rect 26738 35646 26740 35698
rect 26684 35364 26740 35646
rect 26684 35298 26740 35308
rect 26684 34916 26740 34926
rect 26684 34822 26740 34860
rect 26572 33966 26574 34018
rect 26626 33966 26628 34018
rect 26572 32900 26628 33966
rect 26684 34468 26740 34478
rect 26684 33908 26740 34412
rect 26684 33842 26740 33852
rect 26796 33458 26852 36204
rect 26796 33406 26798 33458
rect 26850 33406 26852 33458
rect 26796 33394 26852 33406
rect 26908 33124 26964 36988
rect 27132 36932 27188 39228
rect 27804 38834 27860 40572
rect 27916 40404 27972 40414
rect 27916 40310 27972 40348
rect 27804 38782 27806 38834
rect 27858 38782 27860 38834
rect 27804 38500 27860 38782
rect 28140 38836 28196 38846
rect 28140 38742 28196 38780
rect 28252 38668 28308 43596
rect 28476 41748 28532 47182
rect 28700 46676 28756 46686
rect 28700 46562 28756 46620
rect 28700 46510 28702 46562
rect 28754 46510 28756 46562
rect 28588 45108 28644 45118
rect 28588 45014 28644 45052
rect 28588 44772 28644 44782
rect 28588 44436 28644 44716
rect 28588 43650 28644 44380
rect 28588 43598 28590 43650
rect 28642 43598 28644 43650
rect 28588 43586 28644 43598
rect 27804 38434 27860 38444
rect 28140 38612 28308 38668
rect 28364 41692 28532 41748
rect 28588 42532 28644 42542
rect 28700 42532 28756 46510
rect 28644 42476 28756 42532
rect 28364 39618 28420 41692
rect 28476 41186 28532 41198
rect 28476 41134 28478 41186
rect 28530 41134 28532 41186
rect 28476 40516 28532 41134
rect 28476 40450 28532 40460
rect 28588 39956 28644 42476
rect 28700 41970 28756 41982
rect 28700 41918 28702 41970
rect 28754 41918 28756 41970
rect 28700 41860 28756 41918
rect 28700 41794 28756 41804
rect 28700 41300 28756 41310
rect 28700 40402 28756 41244
rect 28700 40350 28702 40402
rect 28754 40350 28756 40402
rect 28700 40338 28756 40350
rect 28588 39890 28644 39900
rect 28476 39732 28532 39742
rect 28476 39638 28532 39676
rect 28364 39566 28366 39618
rect 28418 39566 28420 39618
rect 27916 38050 27972 38062
rect 27916 37998 27918 38050
rect 27970 37998 27972 38050
rect 27916 37940 27972 37998
rect 27468 37828 27524 37838
rect 27916 37828 27972 37884
rect 27468 37826 27972 37828
rect 27468 37774 27470 37826
rect 27522 37774 27972 37826
rect 27468 37772 27972 37774
rect 27468 37762 27524 37772
rect 27468 37380 27524 37390
rect 27020 36876 27188 36932
rect 27356 36932 27412 36942
rect 27020 35924 27076 36876
rect 27020 35858 27076 35868
rect 27132 36482 27188 36494
rect 27132 36430 27134 36482
rect 27186 36430 27188 36482
rect 27020 34802 27076 34814
rect 27020 34750 27022 34802
rect 27074 34750 27076 34802
rect 27020 34692 27076 34750
rect 27020 34626 27076 34636
rect 27132 33684 27188 36430
rect 27356 35700 27412 36876
rect 27356 35026 27412 35644
rect 27468 35698 27524 37324
rect 27916 36708 27972 37772
rect 28028 37156 28084 37166
rect 28140 37156 28196 38612
rect 28252 38162 28308 38174
rect 28252 38110 28254 38162
rect 28306 38110 28308 38162
rect 28252 37604 28308 38110
rect 28252 37538 28308 37548
rect 28028 37154 28196 37156
rect 28028 37102 28030 37154
rect 28082 37102 28196 37154
rect 28028 37100 28196 37102
rect 28028 37090 28084 37100
rect 27916 36652 28084 36708
rect 27916 36484 27972 36494
rect 27916 36390 27972 36428
rect 27580 36260 27636 36270
rect 27580 35810 27636 36204
rect 27580 35758 27582 35810
rect 27634 35758 27636 35810
rect 27580 35746 27636 35758
rect 27468 35646 27470 35698
rect 27522 35646 27524 35698
rect 27468 35634 27524 35646
rect 27356 34974 27358 35026
rect 27410 34974 27412 35026
rect 27356 34962 27412 34974
rect 27468 35140 27524 35150
rect 27132 33458 27188 33628
rect 27132 33406 27134 33458
rect 27186 33406 27188 33458
rect 27132 33394 27188 33406
rect 26908 33058 26964 33068
rect 26572 32834 26628 32844
rect 25900 32734 25902 32786
rect 25954 32734 25956 32786
rect 25900 32722 25956 32734
rect 25452 32562 25620 32564
rect 25452 32510 25454 32562
rect 25506 32510 25620 32562
rect 25452 32508 25620 32510
rect 25452 32498 25508 32508
rect 27468 31948 27524 35084
rect 27580 33346 27636 33358
rect 27580 33294 27582 33346
rect 27634 33294 27636 33346
rect 27580 33236 27636 33294
rect 27636 33180 27972 33236
rect 27580 33170 27636 33180
rect 27916 32786 27972 33180
rect 27916 32734 27918 32786
rect 27970 32734 27972 32786
rect 27916 32722 27972 32734
rect 26684 31892 27524 31948
rect 25452 31668 25508 31678
rect 25116 31612 25284 31668
rect 24892 31154 24948 31164
rect 25004 31554 25060 31566
rect 25004 31502 25006 31554
rect 25058 31502 25060 31554
rect 25004 31444 25060 31502
rect 25116 31444 25172 31454
rect 25004 31388 25116 31444
rect 22820 30828 22932 30884
rect 23996 30994 24388 30996
rect 23996 30942 24222 30994
rect 24274 30942 24388 30994
rect 23996 30940 24388 30942
rect 22764 30790 22820 30828
rect 21868 30324 21924 30334
rect 21756 30322 21924 30324
rect 21756 30270 21870 30322
rect 21922 30270 21924 30322
rect 21756 30268 21924 30270
rect 21868 30258 21924 30268
rect 23884 30324 23940 30334
rect 23996 30324 24052 30940
rect 24220 30930 24276 30940
rect 24668 30884 24724 30894
rect 24668 30790 24724 30828
rect 24332 30324 24388 30334
rect 23884 30322 24052 30324
rect 23884 30270 23886 30322
rect 23938 30270 24052 30322
rect 23884 30268 24052 30270
rect 24108 30268 24332 30324
rect 23660 30210 23716 30222
rect 23660 30158 23662 30210
rect 23714 30158 23716 30210
rect 22988 30100 23044 30110
rect 22988 30006 23044 30044
rect 23660 30100 23716 30158
rect 23660 30034 23716 30044
rect 20972 29922 21028 29932
rect 23884 29650 23940 30268
rect 23884 29598 23886 29650
rect 23938 29598 23940 29650
rect 23884 29586 23940 29598
rect 20412 28590 20414 28642
rect 20466 28590 20468 28642
rect 20412 28578 20468 28590
rect 20636 29428 20692 29438
rect 20636 28530 20692 29372
rect 22092 29428 22148 29438
rect 22092 29334 22148 29372
rect 22540 29426 22596 29438
rect 22540 29374 22542 29426
rect 22594 29374 22596 29426
rect 22540 29092 22596 29374
rect 24108 29428 24164 30268
rect 24332 30258 24388 30268
rect 24556 30212 24612 30222
rect 24332 30098 24388 30110
rect 24332 30046 24334 30098
rect 24386 30046 24388 30098
rect 24108 29426 24276 29428
rect 24108 29374 24110 29426
rect 24162 29374 24276 29426
rect 24108 29372 24276 29374
rect 24108 29362 24164 29372
rect 22540 29026 22596 29036
rect 23548 29204 23604 29214
rect 20636 28478 20638 28530
rect 20690 28478 20692 28530
rect 20636 28466 20692 28478
rect 23212 28756 23268 28766
rect 23212 28418 23268 28700
rect 23548 28530 23604 29148
rect 23772 29202 23828 29214
rect 23772 29150 23774 29202
rect 23826 29150 23828 29202
rect 23772 28756 23828 29150
rect 24220 28980 24276 29372
rect 24332 29204 24388 30046
rect 24556 30098 24612 30156
rect 25004 30100 25060 31388
rect 25116 31378 25172 31388
rect 25228 31220 25284 31612
rect 25452 31574 25508 31612
rect 25564 31554 25620 31566
rect 25788 31556 25844 31566
rect 25564 31502 25566 31554
rect 25618 31502 25620 31554
rect 25564 31444 25620 31502
rect 25116 31164 25284 31220
rect 25340 31388 25620 31444
rect 25676 31554 25844 31556
rect 25676 31502 25790 31554
rect 25842 31502 25844 31554
rect 25676 31500 25844 31502
rect 25116 30324 25172 31164
rect 25340 30884 25396 31388
rect 25340 30790 25396 30828
rect 25676 30660 25732 31500
rect 25788 31490 25844 31500
rect 26460 31556 26516 31566
rect 26684 31556 26740 31892
rect 28028 31780 28084 36652
rect 28140 36484 28196 37100
rect 28364 36932 28420 39566
rect 28812 38668 28868 48636
rect 28924 48244 28980 48254
rect 28924 48150 28980 48188
rect 28924 48018 28980 48030
rect 28924 47966 28926 48018
rect 28978 47966 28980 48018
rect 28924 45220 28980 47966
rect 29036 46564 29092 46574
rect 29036 46470 29092 46508
rect 29036 45220 29092 45230
rect 28924 45218 29092 45220
rect 28924 45166 29038 45218
rect 29090 45166 29092 45218
rect 28924 45164 29092 45166
rect 29036 45154 29092 45164
rect 29148 44436 29204 49420
rect 29260 49364 29316 49374
rect 29260 49138 29316 49308
rect 29260 49086 29262 49138
rect 29314 49086 29316 49138
rect 29260 49074 29316 49086
rect 29708 48802 29764 49644
rect 29708 48750 29710 48802
rect 29762 48750 29764 48802
rect 29484 48244 29540 48254
rect 29708 48244 29764 48750
rect 29820 48580 29876 49756
rect 30044 49700 30100 49710
rect 29932 49698 30100 49700
rect 29932 49646 30046 49698
rect 30098 49646 30100 49698
rect 29932 49644 30100 49646
rect 29932 49252 29988 49644
rect 30044 49634 30100 49644
rect 29932 49186 29988 49196
rect 30044 49028 30100 49038
rect 30044 48934 30100 48972
rect 29820 48524 30100 48580
rect 29484 48242 29764 48244
rect 29484 48190 29486 48242
rect 29538 48190 29764 48242
rect 29484 48188 29764 48190
rect 29932 48354 29988 48366
rect 29932 48302 29934 48354
rect 29986 48302 29988 48354
rect 29932 48244 29988 48302
rect 29484 48178 29540 48188
rect 29932 48178 29988 48188
rect 29820 48018 29876 48030
rect 29820 47966 29822 48018
rect 29874 47966 29876 48018
rect 29260 47460 29316 47470
rect 29260 47366 29316 47404
rect 29596 47460 29652 47470
rect 29260 45780 29316 45790
rect 29260 45686 29316 45724
rect 29484 45106 29540 45118
rect 29484 45054 29486 45106
rect 29538 45054 29540 45106
rect 29260 44436 29316 44446
rect 29484 44436 29540 45054
rect 29148 44434 29428 44436
rect 29148 44382 29262 44434
rect 29314 44382 29428 44434
rect 29148 44380 29428 44382
rect 29260 44370 29316 44380
rect 29148 43540 29204 43550
rect 29148 43538 29316 43540
rect 29148 43486 29150 43538
rect 29202 43486 29316 43538
rect 29148 43484 29316 43486
rect 29148 43474 29204 43484
rect 29148 42642 29204 42654
rect 29148 42590 29150 42642
rect 29202 42590 29204 42642
rect 29148 41524 29204 42590
rect 29148 40852 29204 41468
rect 29260 42082 29316 43484
rect 29372 42978 29428 44380
rect 29484 44370 29540 44380
rect 29372 42926 29374 42978
rect 29426 42926 29428 42978
rect 29372 42914 29428 42926
rect 29596 42756 29652 47404
rect 29708 46116 29764 46126
rect 29820 46116 29876 47966
rect 29932 47572 29988 47582
rect 29932 47478 29988 47516
rect 30044 46564 30100 48524
rect 30156 48354 30212 49756
rect 30268 49718 30324 49756
rect 30716 49812 30772 49822
rect 30716 49718 30772 49756
rect 30828 49810 30884 49822
rect 30828 49758 30830 49810
rect 30882 49758 30884 49810
rect 30828 49588 30884 49758
rect 30716 49532 30884 49588
rect 30380 49140 30436 49150
rect 30268 49084 30380 49140
rect 30268 48914 30324 49084
rect 30380 49074 30436 49084
rect 30604 49028 30660 49038
rect 30716 49028 30772 49532
rect 30660 48972 30772 49028
rect 30828 49026 30884 49038
rect 30828 48974 30830 49026
rect 30882 48974 30884 49026
rect 30604 48962 30660 48972
rect 30268 48862 30270 48914
rect 30322 48862 30324 48914
rect 30268 48850 30324 48862
rect 30828 48804 30884 48974
rect 30828 48738 30884 48748
rect 30156 48302 30158 48354
rect 30210 48302 30212 48354
rect 30156 48290 30212 48302
rect 30268 48692 30324 48702
rect 30156 47684 30212 47694
rect 30156 47590 30212 47628
rect 30268 47458 30324 48636
rect 30604 48580 30660 48590
rect 30940 48580 30996 51436
rect 31164 51492 31220 51502
rect 31220 51436 31332 51492
rect 31164 51426 31220 51436
rect 31052 51378 31108 51390
rect 31052 51326 31054 51378
rect 31106 51326 31108 51378
rect 31052 50708 31108 51326
rect 31276 51378 31332 51436
rect 31276 51326 31278 51378
rect 31330 51326 31332 51378
rect 31276 51314 31332 51326
rect 31164 51268 31220 51278
rect 31164 51174 31220 51212
rect 31388 51156 31444 51660
rect 31388 51090 31444 51100
rect 31052 50652 31220 50708
rect 31164 50594 31220 50652
rect 31164 50542 31166 50594
rect 31218 50542 31220 50594
rect 31052 50482 31108 50494
rect 31052 50430 31054 50482
rect 31106 50430 31108 50482
rect 31052 50372 31108 50430
rect 31052 50306 31108 50316
rect 31164 49810 31220 50542
rect 31164 49758 31166 49810
rect 31218 49758 31220 49810
rect 30660 48524 30996 48580
rect 30492 48356 30548 48366
rect 30604 48356 30660 48524
rect 30492 48354 30660 48356
rect 30492 48302 30494 48354
rect 30546 48302 30660 48354
rect 30492 48300 30660 48302
rect 30492 48290 30548 48300
rect 30268 47406 30270 47458
rect 30322 47406 30324 47458
rect 30268 47068 30324 47406
rect 30828 48244 30884 48254
rect 30828 47348 30884 48188
rect 30940 47682 30996 48524
rect 30940 47630 30942 47682
rect 30994 47630 30996 47682
rect 30940 47618 30996 47630
rect 31052 49476 31108 49486
rect 30828 47282 30884 47292
rect 30268 47012 30996 47068
rect 30828 46676 30884 46686
rect 30828 46582 30884 46620
rect 30492 46564 30548 46574
rect 30044 46508 30492 46564
rect 29932 46116 29988 46126
rect 29820 46060 29932 46116
rect 29708 45668 29764 46060
rect 29932 46050 29988 46060
rect 30156 45892 30212 45902
rect 30044 45780 30100 45790
rect 29708 45574 29764 45612
rect 29932 45724 30044 45780
rect 29708 44882 29764 44894
rect 29708 44830 29710 44882
rect 29762 44830 29764 44882
rect 29708 44772 29764 44830
rect 29708 44706 29764 44716
rect 29820 44322 29876 44334
rect 29820 44270 29822 44322
rect 29874 44270 29876 44322
rect 29708 44212 29764 44222
rect 29708 43650 29764 44156
rect 29708 43598 29710 43650
rect 29762 43598 29764 43650
rect 29708 43586 29764 43598
rect 29708 42980 29764 42990
rect 29820 42980 29876 44270
rect 29932 44324 29988 45724
rect 30044 45686 30100 45724
rect 30044 45220 30100 45230
rect 30156 45220 30212 45836
rect 30492 45556 30548 46508
rect 30940 45778 30996 47012
rect 30940 45726 30942 45778
rect 30994 45726 30996 45778
rect 30940 45714 30996 45726
rect 30044 45218 30212 45220
rect 30044 45166 30046 45218
rect 30098 45166 30212 45218
rect 30044 45164 30212 45166
rect 30268 45500 30548 45556
rect 30604 45668 30660 45678
rect 30044 45154 30100 45164
rect 30268 45108 30324 45500
rect 29932 44258 29988 44268
rect 30156 45052 30324 45108
rect 30604 45106 30660 45612
rect 30828 45220 30884 45230
rect 31052 45220 31108 49420
rect 31164 48242 31220 49758
rect 31500 50482 31556 50494
rect 31500 50430 31502 50482
rect 31554 50430 31556 50482
rect 31500 50372 31556 50430
rect 31276 49364 31332 49374
rect 31276 49026 31332 49308
rect 31276 48974 31278 49026
rect 31330 48974 31332 49026
rect 31276 48962 31332 48974
rect 31388 48804 31444 48814
rect 31388 48710 31444 48748
rect 31164 48190 31166 48242
rect 31218 48190 31220 48242
rect 31164 47460 31220 48190
rect 31164 47394 31220 47404
rect 31276 48356 31332 48366
rect 31500 48356 31556 50316
rect 31612 49476 31668 55692
rect 33292 55468 33348 56030
rect 33516 55972 33572 55982
rect 33516 55878 33572 55916
rect 33740 55468 33796 56142
rect 32732 55412 33348 55468
rect 33628 55412 33796 55468
rect 33852 56082 33908 56094
rect 33852 56030 33854 56082
rect 33906 56030 33908 56082
rect 31948 54628 32004 54638
rect 31948 54514 32004 54572
rect 31948 54462 31950 54514
rect 32002 54462 32004 54514
rect 31948 54450 32004 54462
rect 31948 53732 32004 53742
rect 31948 52946 32004 53676
rect 31948 52894 31950 52946
rect 32002 52894 32004 52946
rect 31948 52882 32004 52894
rect 31724 52834 31780 52846
rect 31724 52782 31726 52834
rect 31778 52782 31780 52834
rect 31724 52724 31780 52782
rect 32284 52836 32340 52846
rect 32284 52742 32340 52780
rect 31724 50482 31780 52668
rect 31724 50430 31726 50482
rect 31778 50430 31780 50482
rect 31724 50418 31780 50430
rect 31836 50484 31892 50494
rect 31836 50390 31892 50428
rect 31612 49410 31668 49420
rect 31276 48354 31556 48356
rect 31276 48302 31278 48354
rect 31330 48302 31556 48354
rect 31276 48300 31556 48302
rect 31612 49140 31668 49150
rect 31164 47236 31220 47246
rect 31276 47236 31332 48300
rect 31612 47682 31668 49084
rect 32172 48468 32228 48478
rect 32060 48244 32116 48254
rect 32060 48150 32116 48188
rect 31612 47630 31614 47682
rect 31666 47630 31668 47682
rect 31612 47618 31668 47630
rect 31220 47180 31332 47236
rect 31388 47570 31444 47582
rect 31388 47518 31390 47570
rect 31442 47518 31444 47570
rect 31164 47142 31220 47180
rect 31276 47012 31332 47022
rect 31276 46898 31332 46956
rect 31276 46846 31278 46898
rect 31330 46846 31332 46898
rect 31276 46834 31332 46846
rect 31388 46898 31444 47518
rect 31948 47570 32004 47582
rect 31948 47518 31950 47570
rect 32002 47518 32004 47570
rect 31388 46846 31390 46898
rect 31442 46846 31444 46898
rect 31388 46834 31444 46846
rect 31500 47348 31556 47358
rect 31164 46674 31220 46686
rect 31164 46622 31166 46674
rect 31218 46622 31220 46674
rect 31164 46564 31220 46622
rect 31164 46498 31220 46508
rect 31500 46452 31556 47292
rect 31276 46396 31556 46452
rect 30828 45218 31108 45220
rect 30828 45166 30830 45218
rect 30882 45166 31108 45218
rect 30828 45164 31108 45166
rect 31164 45890 31220 45902
rect 31164 45838 31166 45890
rect 31218 45838 31220 45890
rect 31164 45780 31220 45838
rect 30828 45154 30884 45164
rect 30604 45054 30606 45106
rect 30658 45054 30660 45106
rect 29708 42978 29876 42980
rect 29708 42926 29710 42978
rect 29762 42926 29876 42978
rect 29708 42924 29876 42926
rect 29708 42914 29764 42924
rect 29596 42700 29764 42756
rect 29260 42030 29262 42082
rect 29314 42030 29316 42082
rect 29260 41748 29316 42030
rect 29260 41300 29316 41692
rect 29372 41300 29428 41310
rect 29260 41298 29428 41300
rect 29260 41246 29374 41298
rect 29426 41246 29428 41298
rect 29260 41244 29428 41246
rect 29148 40786 29204 40796
rect 29372 40628 29428 41244
rect 29372 40562 29428 40572
rect 29260 40180 29316 40190
rect 29260 39618 29316 40124
rect 29596 40180 29652 40190
rect 29260 39566 29262 39618
rect 29314 39566 29316 39618
rect 29260 39554 29316 39566
rect 29372 39620 29428 39630
rect 29372 39506 29428 39564
rect 29596 39618 29652 40124
rect 29596 39566 29598 39618
rect 29650 39566 29652 39618
rect 29596 39554 29652 39566
rect 29372 39454 29374 39506
rect 29426 39454 29428 39506
rect 29372 39396 29428 39454
rect 29372 39330 29428 39340
rect 29596 39060 29652 39070
rect 29596 38966 29652 39004
rect 29148 38948 29204 38958
rect 29148 38854 29204 38892
rect 28364 36708 28420 36876
rect 28700 38612 28868 38668
rect 28476 36708 28532 36718
rect 28364 36706 28532 36708
rect 28364 36654 28478 36706
rect 28530 36654 28532 36706
rect 28364 36652 28532 36654
rect 28476 36642 28532 36652
rect 28140 36482 28308 36484
rect 28140 36430 28142 36482
rect 28194 36430 28308 36482
rect 28140 36428 28308 36430
rect 28140 36418 28196 36428
rect 28140 35028 28196 35038
rect 28140 34934 28196 34972
rect 28140 33460 28196 33470
rect 28140 33366 28196 33404
rect 28140 33012 28196 33022
rect 28252 33012 28308 36428
rect 28364 35364 28420 35374
rect 28700 35364 28756 38612
rect 29708 38274 29764 42700
rect 29820 40964 29876 40974
rect 29820 40962 29988 40964
rect 29820 40910 29822 40962
rect 29874 40910 29988 40962
rect 29820 40908 29988 40910
rect 29820 40898 29876 40908
rect 29820 40628 29876 40638
rect 29820 40402 29876 40572
rect 29820 40350 29822 40402
rect 29874 40350 29876 40402
rect 29820 40338 29876 40350
rect 29708 38222 29710 38274
rect 29762 38222 29764 38274
rect 29708 38210 29764 38222
rect 29820 39394 29876 39406
rect 29820 39342 29822 39394
rect 29874 39342 29876 39394
rect 29596 38050 29652 38062
rect 29596 37998 29598 38050
rect 29650 37998 29652 38050
rect 29260 37940 29316 37950
rect 29596 37940 29652 37998
rect 29316 37884 29652 37940
rect 29708 37940 29764 37950
rect 29820 37940 29876 39342
rect 29708 37938 29876 37940
rect 29708 37886 29710 37938
rect 29762 37886 29876 37938
rect 29708 37884 29876 37886
rect 29932 38948 29988 40908
rect 30044 38948 30100 38958
rect 29932 38946 30100 38948
rect 29932 38894 30046 38946
rect 30098 38894 30100 38946
rect 29932 38892 30100 38894
rect 29260 37846 29316 37884
rect 29372 37716 29428 37726
rect 29260 37268 29316 37278
rect 29148 37266 29316 37268
rect 29148 37214 29262 37266
rect 29314 37214 29316 37266
rect 29148 37212 29316 37214
rect 29148 36482 29204 37212
rect 29260 37202 29316 37212
rect 29260 36596 29316 36634
rect 29260 36530 29316 36540
rect 29148 36430 29150 36482
rect 29202 36430 29204 36482
rect 29036 35924 29092 35934
rect 29036 35830 29092 35868
rect 28924 35700 28980 35710
rect 28924 35606 28980 35644
rect 28364 34130 28420 35308
rect 28476 35308 28756 35364
rect 28476 35140 28532 35308
rect 28476 35074 28532 35084
rect 28588 35140 28644 35150
rect 29148 35140 29204 36430
rect 29260 36370 29316 36382
rect 29260 36318 29262 36370
rect 29314 36318 29316 36370
rect 29260 35364 29316 36318
rect 29260 35298 29316 35308
rect 28588 35138 29204 35140
rect 28588 35086 28590 35138
rect 28642 35086 29204 35138
rect 28588 35084 29204 35086
rect 28588 35074 28644 35084
rect 29260 35028 29316 35038
rect 29148 34916 29204 34926
rect 28476 34804 28532 34814
rect 28476 34710 28532 34748
rect 28364 34078 28366 34130
rect 28418 34078 28420 34130
rect 28364 33460 28420 34078
rect 28700 34130 28756 34142
rect 28700 34078 28702 34130
rect 28754 34078 28756 34130
rect 28700 33908 28756 34078
rect 29036 34132 29092 34142
rect 29036 34038 29092 34076
rect 28700 33842 28756 33852
rect 28364 33394 28420 33404
rect 28476 33346 28532 33358
rect 28476 33294 28478 33346
rect 28530 33294 28532 33346
rect 28476 33236 28532 33294
rect 28532 33180 28756 33236
rect 28476 33170 28532 33180
rect 28196 32956 28308 33012
rect 28140 32946 28196 32956
rect 28700 32786 28756 33180
rect 29148 33234 29204 34860
rect 29260 34914 29316 34972
rect 29260 34862 29262 34914
rect 29314 34862 29316 34914
rect 29260 34850 29316 34862
rect 29372 33572 29428 37660
rect 29484 34916 29540 34926
rect 29484 34822 29540 34860
rect 29708 34914 29764 37884
rect 29820 37156 29876 37166
rect 29932 37156 29988 38892
rect 30044 38882 30100 38892
rect 30156 38668 30212 45052
rect 30492 44548 30548 44558
rect 30268 43538 30324 43550
rect 30268 43486 30270 43538
rect 30322 43486 30324 43538
rect 30268 42644 30324 43486
rect 30492 43428 30548 44492
rect 30604 44324 30660 45054
rect 30940 44996 30996 45006
rect 30604 44258 30660 44268
rect 30828 44940 30940 44996
rect 30380 42644 30436 42654
rect 30268 42588 30380 42644
rect 30268 41972 30324 41982
rect 30268 41878 30324 41916
rect 30380 41298 30436 42588
rect 30492 42532 30548 43372
rect 30716 43538 30772 43550
rect 30716 43486 30718 43538
rect 30770 43486 30772 43538
rect 30604 42868 30660 42878
rect 30604 42754 30660 42812
rect 30604 42702 30606 42754
rect 30658 42702 30660 42754
rect 30604 42690 30660 42702
rect 30716 42756 30772 43486
rect 30828 42866 30884 44940
rect 30940 44930 30996 44940
rect 31164 44772 31220 45724
rect 31052 44716 31220 44772
rect 30940 44324 30996 44334
rect 30940 43316 30996 44268
rect 31052 43538 31108 44716
rect 31276 44660 31332 46396
rect 31500 46116 31556 46126
rect 31388 44884 31444 44894
rect 31388 44790 31444 44828
rect 31276 44604 31444 44660
rect 31164 44324 31220 44334
rect 31164 44322 31332 44324
rect 31164 44270 31166 44322
rect 31218 44270 31332 44322
rect 31164 44268 31332 44270
rect 31164 44258 31220 44268
rect 31276 43762 31332 44268
rect 31388 43988 31444 44604
rect 31500 44322 31556 46060
rect 31612 45892 31668 45902
rect 31612 45798 31668 45836
rect 31836 45780 31892 45790
rect 31724 45724 31836 45780
rect 31724 45330 31780 45724
rect 31836 45686 31892 45724
rect 31724 45278 31726 45330
rect 31778 45278 31780 45330
rect 31724 45266 31780 45278
rect 31836 45444 31892 45454
rect 31500 44270 31502 44322
rect 31554 44270 31556 44322
rect 31500 44258 31556 44270
rect 31836 44210 31892 45388
rect 31948 44996 32004 47518
rect 32060 47460 32116 47470
rect 32172 47460 32228 48412
rect 32060 47458 32228 47460
rect 32060 47406 32062 47458
rect 32114 47406 32228 47458
rect 32060 47404 32228 47406
rect 32060 47394 32116 47404
rect 32620 47236 32676 47246
rect 32508 46004 32564 46014
rect 32508 45890 32564 45948
rect 32508 45838 32510 45890
rect 32562 45838 32564 45890
rect 32508 45826 32564 45838
rect 32620 45892 32676 47180
rect 32732 46114 32788 55412
rect 33068 55300 33124 55310
rect 33068 55206 33124 55244
rect 32956 55186 33012 55198
rect 32956 55134 32958 55186
rect 33010 55134 33012 55186
rect 32956 53842 33012 55134
rect 33180 54628 33236 54638
rect 33180 54534 33236 54572
rect 32956 53790 32958 53842
rect 33010 53790 33012 53842
rect 32956 52948 33012 53790
rect 32956 52882 33012 52892
rect 33292 53730 33348 53742
rect 33292 53678 33294 53730
rect 33346 53678 33348 53730
rect 33292 53620 33348 53678
rect 33292 52164 33348 53564
rect 33404 53620 33460 53630
rect 33628 53620 33684 55412
rect 33740 55298 33796 55310
rect 33740 55246 33742 55298
rect 33794 55246 33796 55298
rect 33740 54964 33796 55246
rect 33852 55188 33908 56030
rect 48188 56082 48244 56094
rect 48188 56030 48190 56082
rect 48242 56030 48244 56082
rect 34748 55970 34804 55982
rect 34748 55918 34750 55970
rect 34802 55918 34804 55970
rect 34076 55300 34132 55310
rect 34076 55206 34132 55244
rect 33852 55122 33908 55132
rect 34524 55188 34580 55198
rect 34748 55188 34804 55918
rect 34524 55186 34804 55188
rect 34524 55134 34526 55186
rect 34578 55134 34804 55186
rect 34524 55132 34804 55134
rect 34860 55972 34916 55982
rect 33740 54908 34244 54964
rect 33852 54740 33908 54750
rect 33852 54292 33908 54684
rect 34188 54628 34244 54908
rect 34524 54628 34580 55132
rect 34860 54628 34916 55916
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 48188 55522 48244 56030
rect 48188 55470 48190 55522
rect 48242 55470 48244 55522
rect 48188 55458 48244 55470
rect 48412 55412 48468 59200
rect 48972 56308 49028 56318
rect 49084 56308 49140 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49196 56308 49252 56318
rect 49084 56252 49196 56308
rect 48972 56214 49028 56252
rect 49196 56242 49252 56252
rect 48412 55346 48468 55356
rect 49532 56084 49588 56094
rect 34188 54626 34580 54628
rect 34188 54574 34190 54626
rect 34242 54574 34580 54626
rect 34188 54572 34580 54574
rect 34636 54572 34916 54628
rect 35084 55298 35140 55310
rect 35084 55246 35086 55298
rect 35138 55246 35140 55298
rect 34076 54514 34132 54526
rect 34076 54462 34078 54514
rect 34130 54462 34132 54514
rect 34076 54404 34132 54462
rect 34076 54338 34132 54348
rect 33852 53730 33908 54236
rect 33852 53678 33854 53730
rect 33906 53678 33908 53730
rect 33852 53666 33908 53678
rect 33404 53618 33684 53620
rect 33404 53566 33406 53618
rect 33458 53566 33684 53618
rect 33404 53564 33684 53566
rect 33404 53554 33460 53564
rect 33628 53170 33684 53564
rect 34188 53618 34244 54572
rect 34636 53842 34692 54572
rect 34636 53790 34638 53842
rect 34690 53790 34692 53842
rect 34636 53778 34692 53790
rect 34412 53732 34468 53742
rect 34412 53638 34468 53676
rect 34972 53730 35028 53742
rect 34972 53678 34974 53730
rect 35026 53678 35028 53730
rect 34188 53566 34190 53618
rect 34242 53566 34244 53618
rect 34188 53554 34244 53566
rect 33628 53118 33630 53170
rect 33682 53118 33684 53170
rect 33628 53106 33684 53118
rect 33404 52948 33460 52958
rect 33740 52948 33796 52958
rect 33404 52946 33796 52948
rect 33404 52894 33406 52946
rect 33458 52894 33742 52946
rect 33794 52894 33796 52946
rect 33404 52892 33796 52894
rect 33404 52882 33460 52892
rect 33292 52108 33684 52164
rect 33180 51156 33236 51166
rect 32956 50484 33012 50494
rect 32956 50390 33012 50428
rect 33068 50482 33124 50494
rect 33068 50430 33070 50482
rect 33122 50430 33124 50482
rect 32732 46062 32734 46114
rect 32786 46062 32788 46114
rect 32732 46050 32788 46062
rect 33068 48804 33124 50430
rect 33180 49026 33236 51100
rect 33292 50596 33348 50606
rect 33292 50502 33348 50540
rect 33628 49252 33684 52108
rect 33516 49196 33684 49252
rect 33180 48974 33182 49026
rect 33234 48974 33236 49026
rect 33180 48962 33236 48974
rect 33292 49028 33348 49038
rect 32844 45892 32900 45902
rect 32620 45836 32788 45892
rect 31948 44930 32004 44940
rect 32284 44994 32340 45006
rect 32284 44942 32286 44994
rect 32338 44942 32340 44994
rect 32284 44324 32340 44942
rect 32284 44258 32340 44268
rect 31836 44158 31838 44210
rect 31890 44158 31892 44210
rect 31836 44146 31892 44158
rect 31388 43932 31892 43988
rect 31276 43710 31278 43762
rect 31330 43710 31332 43762
rect 31276 43698 31332 43710
rect 31052 43486 31054 43538
rect 31106 43486 31108 43538
rect 31052 43474 31108 43486
rect 30940 43260 31108 43316
rect 30828 42814 30830 42866
rect 30882 42814 30884 42866
rect 30828 42802 30884 42814
rect 30716 42690 30772 42700
rect 30828 42532 30884 42542
rect 30492 42530 30884 42532
rect 30492 42478 30830 42530
rect 30882 42478 30884 42530
rect 30492 42476 30884 42478
rect 30380 41246 30382 41298
rect 30434 41246 30436 41298
rect 30380 41234 30436 41246
rect 30492 41074 30548 41086
rect 30492 41022 30494 41074
rect 30546 41022 30548 41074
rect 30268 40962 30324 40974
rect 30268 40910 30270 40962
rect 30322 40910 30324 40962
rect 30268 39956 30324 40910
rect 30268 39890 30324 39900
rect 30492 40068 30548 41022
rect 30828 41074 30884 42476
rect 30940 42530 30996 42542
rect 30940 42478 30942 42530
rect 30994 42478 30996 42530
rect 30940 42084 30996 42478
rect 30940 41412 30996 42028
rect 31052 41524 31108 43260
rect 31724 42866 31780 42878
rect 31724 42814 31726 42866
rect 31778 42814 31780 42866
rect 31388 42644 31444 42654
rect 31388 42550 31444 42588
rect 31612 42532 31668 42542
rect 31612 42438 31668 42476
rect 31500 42196 31556 42206
rect 31500 42194 31668 42196
rect 31500 42142 31502 42194
rect 31554 42142 31668 42194
rect 31500 42140 31668 42142
rect 31500 42130 31556 42140
rect 31052 41468 31220 41524
rect 30940 41356 31108 41412
rect 31052 41186 31108 41356
rect 31052 41134 31054 41186
rect 31106 41134 31108 41186
rect 31052 41122 31108 41134
rect 30828 41022 30830 41074
rect 30882 41022 30884 41074
rect 30828 40180 30884 41022
rect 30940 40852 30996 40862
rect 30940 40402 30996 40796
rect 30940 40350 30942 40402
rect 30994 40350 30996 40402
rect 30940 40338 30996 40350
rect 31052 40180 31108 40190
rect 30828 40124 31052 40180
rect 31052 40114 31108 40124
rect 29820 37154 29988 37156
rect 29820 37102 29822 37154
rect 29874 37102 29988 37154
rect 29820 37100 29988 37102
rect 30044 38612 30212 38668
rect 30268 39620 30324 39630
rect 30268 38722 30324 39564
rect 30380 39618 30436 39630
rect 30380 39566 30382 39618
rect 30434 39566 30436 39618
rect 30380 39396 30436 39566
rect 30380 39330 30436 39340
rect 30268 38670 30270 38722
rect 30322 38670 30324 38722
rect 30268 38658 30324 38670
rect 29820 37044 29876 37100
rect 29820 36978 29876 36988
rect 30044 35700 30100 38612
rect 30268 37156 30324 37166
rect 30268 37062 30324 37100
rect 30268 36596 30324 36606
rect 30492 36596 30548 40012
rect 30716 40012 30996 40068
rect 30604 38948 30660 38958
rect 30604 38834 30660 38892
rect 30604 38782 30606 38834
rect 30658 38782 30660 38834
rect 30604 38770 30660 38782
rect 30716 38052 30772 40012
rect 30940 39956 30996 40012
rect 31164 39956 31220 41468
rect 31500 41074 31556 41086
rect 31500 41022 31502 41074
rect 31554 41022 31556 41074
rect 31500 40628 31556 41022
rect 31612 40964 31668 42140
rect 31724 42082 31780 42814
rect 31724 42030 31726 42082
rect 31778 42030 31780 42082
rect 31724 42018 31780 42030
rect 31612 40898 31668 40908
rect 31500 40562 31556 40572
rect 31836 40404 31892 43932
rect 32284 43540 32340 43550
rect 32284 43446 32340 43484
rect 31948 43428 32004 43438
rect 31948 43334 32004 43372
rect 32620 43428 32676 43438
rect 32620 42866 32676 43372
rect 32620 42814 32622 42866
rect 32674 42814 32676 42866
rect 32620 42802 32676 42814
rect 32172 42530 32228 42542
rect 32172 42478 32174 42530
rect 32226 42478 32228 42530
rect 32172 42420 32228 42478
rect 32228 42364 32452 42420
rect 32172 42354 32228 42364
rect 32172 41970 32228 41982
rect 32172 41918 32174 41970
rect 32226 41918 32228 41970
rect 32172 41412 32228 41918
rect 32172 41346 32228 41356
rect 32396 41300 32452 42364
rect 32396 41206 32452 41244
rect 32508 41860 32564 41870
rect 32172 41186 32228 41198
rect 32172 41134 32174 41186
rect 32226 41134 32228 41186
rect 32172 40628 32228 41134
rect 32172 40562 32228 40572
rect 32508 41186 32564 41804
rect 32508 41134 32510 41186
rect 32562 41134 32564 41186
rect 30940 39900 31220 39956
rect 31500 40348 31892 40404
rect 32284 40402 32340 40414
rect 32284 40350 32286 40402
rect 32338 40350 32340 40402
rect 30828 39844 30884 39854
rect 30828 39732 30884 39788
rect 30828 39730 31108 39732
rect 30828 39678 30830 39730
rect 30882 39678 31108 39730
rect 30828 39676 31108 39678
rect 30828 39666 30884 39676
rect 31052 39284 31108 39676
rect 31164 39618 31220 39630
rect 31164 39566 31166 39618
rect 31218 39566 31220 39618
rect 31164 39508 31220 39566
rect 31388 39620 31444 39630
rect 31388 39526 31444 39564
rect 31164 39442 31220 39452
rect 31388 39284 31444 39294
rect 31052 39228 31332 39284
rect 31164 39060 31220 39070
rect 30940 39058 31220 39060
rect 30940 39006 31166 39058
rect 31218 39006 31220 39058
rect 30940 39004 31220 39006
rect 30940 38948 30996 39004
rect 31164 38994 31220 39004
rect 31276 39058 31332 39228
rect 31276 39006 31278 39058
rect 31330 39006 31332 39058
rect 31276 38994 31332 39006
rect 30940 38882 30996 38892
rect 30604 37996 30772 38052
rect 30828 38836 30884 38846
rect 30604 36708 30660 37996
rect 30716 37828 30772 37838
rect 30828 37828 30884 38780
rect 31052 38836 31108 38846
rect 31388 38836 31444 39228
rect 31052 38834 31444 38836
rect 31052 38782 31054 38834
rect 31106 38782 31444 38834
rect 31052 38780 31444 38782
rect 31052 38164 31108 38780
rect 31500 38668 31556 40348
rect 31612 40180 31668 40190
rect 31836 40180 31892 40190
rect 31668 40124 31780 40180
rect 31612 40114 31668 40124
rect 31612 39956 31668 39966
rect 31612 38836 31668 39900
rect 31612 38742 31668 38780
rect 31388 38612 31556 38668
rect 31164 38164 31220 38174
rect 31052 38162 31220 38164
rect 31052 38110 31166 38162
rect 31218 38110 31220 38162
rect 31052 38108 31220 38110
rect 31164 38098 31220 38108
rect 30716 37826 30884 37828
rect 30716 37774 30718 37826
rect 30770 37774 30884 37826
rect 30716 37772 30884 37774
rect 30716 37716 30772 37772
rect 30716 37650 30772 37660
rect 31388 37492 31444 38612
rect 31500 38276 31556 38286
rect 31724 38276 31780 40124
rect 31836 40086 31892 40124
rect 32284 38388 32340 40350
rect 32172 38332 32340 38388
rect 31724 38220 32116 38276
rect 31500 37828 31556 38220
rect 31612 38164 31668 38174
rect 31612 38050 31668 38108
rect 31612 37998 31614 38050
rect 31666 37998 31668 38050
rect 31612 37986 31668 37998
rect 31948 37940 32004 37950
rect 31948 37846 32004 37884
rect 31724 37828 31780 37838
rect 31500 37826 31780 37828
rect 31500 37774 31726 37826
rect 31778 37774 31780 37826
rect 31500 37772 31780 37774
rect 31724 37762 31780 37772
rect 31164 37436 31444 37492
rect 31052 37268 31108 37278
rect 30940 37266 31108 37268
rect 30940 37214 31054 37266
rect 31106 37214 31108 37266
rect 30940 37212 31108 37214
rect 30716 37156 30772 37166
rect 30716 37062 30772 37100
rect 30604 36652 30772 36708
rect 30156 36594 30548 36596
rect 30156 36542 30270 36594
rect 30322 36542 30548 36594
rect 30156 36540 30548 36542
rect 30156 36484 30212 36540
rect 30268 36530 30324 36540
rect 30604 36484 30660 36494
rect 30156 35810 30212 36428
rect 30492 36482 30660 36484
rect 30492 36430 30606 36482
rect 30658 36430 30660 36482
rect 30492 36428 30660 36430
rect 30156 35758 30158 35810
rect 30210 35758 30212 35810
rect 30156 35746 30212 35758
rect 30268 36036 30324 36046
rect 29932 35644 30100 35700
rect 29820 35588 29876 35598
rect 29820 35138 29876 35532
rect 29820 35086 29822 35138
rect 29874 35086 29876 35138
rect 29820 35074 29876 35086
rect 29708 34862 29710 34914
rect 29762 34862 29764 34914
rect 29148 33182 29150 33234
rect 29202 33182 29204 33234
rect 29148 33170 29204 33182
rect 29260 33516 29428 33572
rect 28700 32734 28702 32786
rect 28754 32734 28756 32786
rect 28700 31948 28756 32734
rect 29036 32788 29092 32798
rect 29260 32788 29316 33516
rect 29036 32786 29316 32788
rect 29036 32734 29038 32786
rect 29090 32734 29316 32786
rect 29036 32732 29316 32734
rect 29372 33346 29428 33358
rect 29372 33294 29374 33346
rect 29426 33294 29428 33346
rect 29372 32788 29428 33294
rect 29708 33124 29764 34862
rect 29820 34020 29876 34030
rect 29820 33458 29876 33964
rect 29820 33406 29822 33458
rect 29874 33406 29876 33458
rect 29820 33394 29876 33406
rect 29708 33058 29764 33068
rect 29708 32788 29764 32798
rect 29372 32786 29764 32788
rect 29372 32734 29374 32786
rect 29426 32734 29710 32786
rect 29762 32734 29764 32786
rect 29372 32732 29764 32734
rect 29036 32722 29092 32732
rect 29372 32722 29428 32732
rect 29708 32722 29764 32732
rect 29820 32452 29876 32462
rect 29484 32450 29876 32452
rect 29484 32398 29822 32450
rect 29874 32398 29876 32450
rect 29484 32396 29876 32398
rect 29484 31948 29540 32396
rect 29820 32386 29876 32396
rect 29932 31948 29988 35644
rect 30044 35476 30100 35486
rect 30044 33906 30100 35420
rect 30268 35026 30324 35980
rect 30268 34974 30270 35026
rect 30322 34974 30324 35026
rect 30268 34962 30324 34974
rect 30492 34916 30548 36428
rect 30604 36418 30660 36428
rect 30604 36260 30660 36270
rect 30604 35922 30660 36204
rect 30604 35870 30606 35922
rect 30658 35870 30660 35922
rect 30604 35858 30660 35870
rect 30604 35588 30660 35598
rect 30604 35494 30660 35532
rect 30604 34916 30660 34926
rect 30044 33854 30046 33906
rect 30098 33854 30100 33906
rect 30044 33842 30100 33854
rect 30380 34914 30660 34916
rect 30380 34862 30606 34914
rect 30658 34862 30660 34914
rect 30380 34860 30660 34862
rect 30380 34804 30436 34860
rect 30604 34850 30660 34860
rect 30380 33348 30436 34748
rect 30716 34580 30772 36652
rect 30940 36484 30996 37212
rect 31052 37202 31108 37212
rect 30940 36260 30996 36428
rect 31052 36932 31108 36942
rect 31052 36482 31108 36876
rect 31052 36430 31054 36482
rect 31106 36430 31108 36482
rect 31052 36418 31108 36430
rect 30940 36194 30996 36204
rect 30940 36036 30996 36046
rect 30940 35698 30996 35980
rect 30940 35646 30942 35698
rect 30994 35646 30996 35698
rect 30940 35634 30996 35646
rect 31164 35138 31220 37436
rect 31276 37266 31332 37278
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 35252 31332 37214
rect 31500 37266 31556 37278
rect 31500 37214 31502 37266
rect 31554 37214 31556 37266
rect 31388 37154 31444 37166
rect 31388 37102 31390 37154
rect 31442 37102 31444 37154
rect 31388 35700 31444 37102
rect 31500 36932 31556 37214
rect 31612 37266 31668 37278
rect 31612 37214 31614 37266
rect 31666 37214 31668 37266
rect 31612 37156 31668 37214
rect 31612 37090 31668 37100
rect 31500 36866 31556 36876
rect 32060 36036 32116 38220
rect 32172 36820 32228 38332
rect 32284 38164 32340 38174
rect 32284 38070 32340 38108
rect 32172 36754 32228 36764
rect 32396 37156 32452 37166
rect 32396 36482 32452 37100
rect 32396 36430 32398 36482
rect 32450 36430 32452 36482
rect 32396 36418 32452 36430
rect 32508 36372 32564 41134
rect 32620 38052 32676 38062
rect 32620 37958 32676 37996
rect 32732 37828 32788 45836
rect 32844 45444 32900 45836
rect 32844 45378 32900 45388
rect 33068 41074 33124 48748
rect 33292 48802 33348 48972
rect 33292 48750 33294 48802
rect 33346 48750 33348 48802
rect 33292 48738 33348 48750
rect 33404 49026 33460 49038
rect 33404 48974 33406 49026
rect 33458 48974 33460 49026
rect 33404 47684 33460 48974
rect 33516 48804 33572 49196
rect 33628 49026 33684 49038
rect 33628 48974 33630 49026
rect 33682 48974 33684 49026
rect 33628 48916 33684 48974
rect 33740 49028 33796 52892
rect 34188 52946 34244 52958
rect 34188 52894 34190 52946
rect 34242 52894 34244 52946
rect 34076 52836 34132 52846
rect 34076 52162 34132 52780
rect 34188 52274 34244 52894
rect 34188 52222 34190 52274
rect 34242 52222 34244 52274
rect 34188 52210 34244 52222
rect 34300 52948 34356 52958
rect 34076 52110 34078 52162
rect 34130 52110 34132 52162
rect 34076 52098 34132 52110
rect 34300 52162 34356 52892
rect 34748 52948 34804 52958
rect 34972 52948 35028 53678
rect 35084 53620 35140 55246
rect 35420 55298 35476 55310
rect 35420 55246 35422 55298
rect 35474 55246 35476 55298
rect 35196 54402 35252 54414
rect 35196 54350 35198 54402
rect 35250 54350 35252 54402
rect 35196 54292 35252 54350
rect 35420 54404 35476 55246
rect 36988 55300 37044 55310
rect 36988 55206 37044 55244
rect 37212 55298 37268 55310
rect 37212 55246 37214 55298
rect 37266 55246 37268 55298
rect 35532 55076 35588 55086
rect 35532 55074 35700 55076
rect 35532 55022 35534 55074
rect 35586 55022 35700 55074
rect 35532 55020 35700 55022
rect 35532 55010 35588 55020
rect 35644 54514 35700 55020
rect 37212 54516 37268 55246
rect 39004 55298 39060 55310
rect 39004 55246 39006 55298
rect 39058 55246 39060 55298
rect 35644 54462 35646 54514
rect 35698 54462 35700 54514
rect 35644 54450 35700 54462
rect 37100 54514 37268 54516
rect 37100 54462 37214 54514
rect 37266 54462 37268 54514
rect 37100 54460 37268 54462
rect 35420 54338 35476 54348
rect 35196 54226 35252 54236
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 36092 53842 36148 53854
rect 36092 53790 36094 53842
rect 36146 53790 36148 53842
rect 35084 53554 35140 53564
rect 35868 53730 35924 53742
rect 35868 53678 35870 53730
rect 35922 53678 35924 53730
rect 35868 53620 35924 53678
rect 36092 53732 36148 53790
rect 36092 53666 36148 53676
rect 34748 52854 34804 52892
rect 34860 52892 34972 52948
rect 34636 52836 34692 52846
rect 34636 52742 34692 52780
rect 34860 52612 34916 52892
rect 34972 52882 35028 52892
rect 34300 52110 34302 52162
rect 34354 52110 34356 52162
rect 34300 51378 34356 52110
rect 34636 52556 34916 52612
rect 35084 52722 35140 52734
rect 35084 52670 35086 52722
rect 35138 52670 35140 52722
rect 34636 52162 34692 52556
rect 34636 52110 34638 52162
rect 34690 52110 34692 52162
rect 34636 52098 34692 52110
rect 34860 52388 34916 52398
rect 34300 51326 34302 51378
rect 34354 51326 34356 51378
rect 34300 51314 34356 51326
rect 34076 51268 34132 51278
rect 34076 51174 34132 51212
rect 34748 51156 34804 51166
rect 34748 51062 34804 51100
rect 34860 50818 34916 52332
rect 35084 52164 35140 52670
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35084 52098 35140 52108
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 34860 50766 34862 50818
rect 34914 50766 34916 50818
rect 34860 50754 34916 50766
rect 33964 50596 34020 50606
rect 34524 50596 34580 50606
rect 33964 50502 34020 50540
rect 34412 50594 34580 50596
rect 34412 50542 34526 50594
rect 34578 50542 34580 50594
rect 34412 50540 34580 50542
rect 33852 50482 33908 50494
rect 33852 50430 33854 50482
rect 33906 50430 33908 50482
rect 33852 49812 33908 50430
rect 34412 50428 34468 50540
rect 34524 50530 34580 50540
rect 34188 50372 34468 50428
rect 34188 50034 34244 50372
rect 34188 49982 34190 50034
rect 34242 49982 34244 50034
rect 34188 49970 34244 49982
rect 35420 50036 35476 50046
rect 35420 49942 35476 49980
rect 35532 49922 35588 49934
rect 35532 49870 35534 49922
rect 35586 49870 35588 49922
rect 34412 49812 34468 49822
rect 33852 49810 34468 49812
rect 33852 49758 34414 49810
rect 34466 49758 34468 49810
rect 33852 49756 34468 49758
rect 35532 49812 35588 49870
rect 35644 49812 35700 49822
rect 35532 49756 35644 49812
rect 34076 49588 34132 49598
rect 34076 49586 34244 49588
rect 34076 49534 34078 49586
rect 34130 49534 34244 49586
rect 34076 49532 34244 49534
rect 34076 49522 34132 49532
rect 34076 49028 34132 49038
rect 33740 48972 34020 49028
rect 33628 48860 33908 48916
rect 33516 48748 33684 48804
rect 33628 48020 33684 48748
rect 33852 48244 33908 48860
rect 33852 48178 33908 48188
rect 33964 48020 34020 48972
rect 34076 48934 34132 48972
rect 34188 48466 34244 49532
rect 34412 49364 34468 49756
rect 35644 49746 35700 49756
rect 35756 49810 35812 49822
rect 35756 49758 35758 49810
rect 35810 49758 35812 49810
rect 35420 49700 35476 49710
rect 35420 49586 35476 49644
rect 35420 49534 35422 49586
rect 35474 49534 35476 49586
rect 35420 49522 35476 49534
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 34412 49308 34692 49364
rect 35196 49354 35460 49364
rect 34524 49140 34580 49150
rect 34524 49026 34580 49084
rect 34524 48974 34526 49026
rect 34578 48974 34580 49026
rect 34524 48962 34580 48974
rect 34636 49028 34692 49308
rect 34972 49028 35028 49038
rect 34636 49026 35028 49028
rect 34636 48974 34974 49026
rect 35026 48974 35028 49026
rect 34636 48972 35028 48974
rect 34188 48414 34190 48466
rect 34242 48414 34244 48466
rect 34188 48402 34244 48414
rect 34076 48354 34132 48366
rect 34076 48302 34078 48354
rect 34130 48302 34132 48354
rect 34076 48244 34132 48302
rect 34076 48178 34132 48188
rect 33628 47964 33908 48020
rect 33964 47964 34132 48020
rect 33404 47618 33460 47628
rect 33628 47796 33684 47806
rect 33516 45892 33572 45902
rect 33516 45798 33572 45836
rect 33628 43652 33684 47740
rect 33740 45780 33796 45790
rect 33740 45686 33796 45724
rect 33852 45668 33908 47964
rect 33964 45668 34020 45678
rect 33852 45666 34020 45668
rect 33852 45614 33966 45666
rect 34018 45614 34020 45666
rect 33852 45612 34020 45614
rect 33964 45602 34020 45612
rect 34076 44772 34132 47964
rect 34300 48018 34356 48030
rect 34300 47966 34302 48018
rect 34354 47966 34356 48018
rect 34300 47684 34356 47966
rect 34300 47618 34356 47628
rect 34972 46788 35028 48972
rect 35420 49026 35476 49038
rect 35420 48974 35422 49026
rect 35474 48974 35476 49026
rect 35420 48468 35476 48974
rect 35420 48402 35476 48412
rect 35532 49028 35588 49038
rect 35532 48354 35588 48972
rect 35756 49026 35812 49758
rect 35868 49250 35924 53564
rect 36428 53508 36484 53518
rect 36428 53414 36484 53452
rect 36316 52948 36372 52958
rect 36316 52834 36372 52892
rect 36764 52948 36820 52958
rect 37100 52948 37156 54460
rect 37212 54450 37268 54460
rect 37772 55186 37828 55198
rect 37772 55134 37774 55186
rect 37826 55134 37828 55186
rect 37772 54404 37828 55134
rect 37772 54338 37828 54348
rect 38108 54514 38164 54526
rect 38108 54462 38110 54514
rect 38162 54462 38164 54514
rect 37324 53842 37380 53854
rect 37324 53790 37326 53842
rect 37378 53790 37380 53842
rect 37212 53730 37268 53742
rect 37212 53678 37214 53730
rect 37266 53678 37268 53730
rect 37212 53620 37268 53678
rect 37324 53732 37380 53790
rect 37996 53844 38052 53854
rect 37996 53750 38052 53788
rect 37324 53666 37380 53676
rect 37212 53554 37268 53564
rect 38108 53620 38164 54462
rect 38444 54404 38500 54414
rect 38444 54310 38500 54348
rect 36764 52946 36932 52948
rect 36764 52894 36766 52946
rect 36818 52894 36932 52946
rect 36764 52892 36932 52894
rect 36764 52882 36820 52892
rect 36316 52782 36318 52834
rect 36370 52782 36372 52834
rect 36316 52770 36372 52782
rect 36092 51380 36148 51390
rect 36092 51286 36148 51324
rect 36428 51378 36484 51390
rect 36428 51326 36430 51378
rect 36482 51326 36484 51378
rect 35868 49198 35870 49250
rect 35922 49198 35924 49250
rect 35868 49186 35924 49198
rect 36428 49812 36484 51326
rect 36876 50484 36932 52892
rect 37100 52882 37156 52892
rect 38108 52388 38164 53564
rect 38668 54290 38724 54302
rect 38668 54238 38670 54290
rect 38722 54238 38724 54290
rect 38668 53060 38724 54238
rect 38780 53730 38836 53742
rect 38780 53678 38782 53730
rect 38834 53678 38836 53730
rect 38780 53284 38836 53678
rect 38780 53228 38948 53284
rect 38892 53170 38948 53228
rect 38892 53118 38894 53170
rect 38946 53118 38948 53170
rect 38892 53106 38948 53118
rect 39004 53172 39060 55246
rect 39564 55298 39620 55310
rect 40236 55300 40292 55310
rect 39564 55246 39566 55298
rect 39618 55246 39620 55298
rect 39452 53620 39508 53630
rect 39564 53620 39620 55246
rect 39900 55298 40292 55300
rect 39900 55246 40238 55298
rect 40290 55246 40292 55298
rect 39900 55244 40292 55246
rect 39900 54404 39956 55244
rect 40236 55234 40292 55244
rect 48748 55298 48804 55310
rect 48748 55246 48750 55298
rect 48802 55246 48804 55298
rect 41020 55188 41076 55198
rect 41020 55094 41076 55132
rect 42476 55188 42532 55198
rect 42028 55074 42084 55086
rect 42028 55022 42030 55074
rect 42082 55022 42084 55074
rect 41580 54514 41636 54526
rect 41580 54462 41582 54514
rect 41634 54462 41636 54514
rect 39788 53956 39844 53966
rect 39788 53842 39844 53900
rect 39788 53790 39790 53842
rect 39842 53790 39844 53842
rect 39788 53778 39844 53790
rect 39900 53730 39956 54348
rect 41356 54402 41412 54414
rect 41356 54350 41358 54402
rect 41410 54350 41412 54402
rect 41356 53844 41412 54350
rect 41356 53750 41412 53788
rect 39900 53678 39902 53730
rect 39954 53678 39956 53730
rect 39900 53666 39956 53678
rect 39508 53564 39620 53620
rect 39452 53526 39508 53564
rect 41580 53506 41636 54462
rect 42028 54180 42084 55022
rect 42140 55076 42196 55086
rect 42140 54982 42196 55020
rect 42252 55076 42308 55086
rect 42252 55074 42420 55076
rect 42252 55022 42254 55074
rect 42306 55022 42420 55074
rect 42252 55020 42420 55022
rect 42252 55010 42308 55020
rect 42252 54516 42308 54526
rect 42252 54422 42308 54460
rect 41692 54124 42308 54180
rect 41692 53954 41748 54124
rect 41692 53902 41694 53954
rect 41746 53902 41748 53954
rect 41692 53890 41748 53902
rect 42252 53954 42308 54124
rect 42252 53902 42254 53954
rect 42306 53902 42308 53954
rect 42252 53890 42308 53902
rect 41580 53454 41582 53506
rect 41634 53454 41636 53506
rect 39004 53170 40068 53172
rect 39004 53118 39006 53170
rect 39058 53118 40068 53170
rect 39004 53116 40068 53118
rect 39004 53106 39060 53116
rect 38780 53060 38836 53070
rect 38668 53058 38836 53060
rect 38668 53006 38782 53058
rect 38834 53006 38836 53058
rect 38668 53004 38836 53006
rect 38780 52994 38836 53004
rect 38108 52322 38164 52332
rect 38444 52724 38500 52734
rect 38444 52162 38500 52668
rect 40012 52274 40068 53116
rect 40012 52222 40014 52274
rect 40066 52222 40068 52274
rect 40012 52210 40068 52222
rect 40908 52276 40964 52286
rect 41580 52276 41636 53454
rect 42028 53732 42084 53742
rect 42364 53732 42420 55020
rect 42476 53954 42532 55132
rect 42924 55188 42980 55198
rect 42476 53902 42478 53954
rect 42530 53902 42532 53954
rect 42476 53890 42532 53902
rect 42588 54292 42644 54302
rect 42028 53730 42420 53732
rect 42028 53678 42030 53730
rect 42082 53678 42420 53730
rect 42028 53676 42420 53678
rect 42028 53508 42084 53676
rect 42028 53442 42084 53452
rect 40908 52274 41636 52276
rect 40908 52222 40910 52274
rect 40962 52222 41636 52274
rect 40908 52220 41636 52222
rect 40908 52210 40964 52220
rect 39116 52164 39172 52174
rect 38444 52110 38446 52162
rect 38498 52110 38500 52162
rect 38444 52098 38500 52110
rect 39004 52162 39172 52164
rect 39004 52110 39118 52162
rect 39170 52110 39172 52162
rect 39004 52108 39172 52110
rect 38556 52050 38612 52062
rect 38556 51998 38558 52050
rect 38610 51998 38612 52050
rect 37548 51940 37604 51950
rect 36988 51492 37044 51502
rect 36988 51398 37044 51436
rect 37548 51490 37604 51884
rect 37548 51438 37550 51490
rect 37602 51438 37604 51490
rect 37548 50596 37604 51438
rect 38332 51490 38388 51502
rect 38332 51438 38334 51490
rect 38386 51438 38388 51490
rect 37884 51380 37940 51390
rect 38332 51380 38388 51438
rect 37884 51378 38388 51380
rect 37884 51326 37886 51378
rect 37938 51326 38388 51378
rect 37884 51324 38388 51326
rect 37884 51314 37940 51324
rect 37548 50530 37604 50540
rect 37660 51156 37716 51166
rect 36876 50428 37380 50484
rect 36876 50260 36932 50270
rect 36876 49922 36932 50204
rect 36876 49870 36878 49922
rect 36930 49870 36932 49922
rect 36876 49858 36932 49870
rect 36428 49698 36484 49756
rect 36428 49646 36430 49698
rect 36482 49646 36484 49698
rect 35756 48974 35758 49026
rect 35810 48974 35812 49026
rect 35644 48804 35700 48814
rect 35644 48466 35700 48748
rect 35644 48414 35646 48466
rect 35698 48414 35700 48466
rect 35644 48402 35700 48414
rect 35756 48468 35812 48974
rect 35868 48468 35924 48478
rect 35756 48466 35924 48468
rect 35756 48414 35870 48466
rect 35922 48414 35924 48466
rect 35756 48412 35924 48414
rect 35868 48402 35924 48412
rect 35532 48302 35534 48354
rect 35586 48302 35588 48354
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35420 46900 35476 46910
rect 35532 46900 35588 48302
rect 36428 48354 36484 49646
rect 36540 49810 36596 49822
rect 36540 49758 36542 49810
rect 36594 49758 36596 49810
rect 36540 48804 36596 49758
rect 36540 48738 36596 48748
rect 36428 48302 36430 48354
rect 36482 48302 36484 48354
rect 36428 48290 36484 48302
rect 36316 48242 36372 48254
rect 36316 48190 36318 48242
rect 36370 48190 36372 48242
rect 36316 47684 36372 48190
rect 36540 48244 36596 48254
rect 37212 48244 37268 48254
rect 36540 47684 36596 48188
rect 36316 47618 36372 47628
rect 36428 47628 36596 47684
rect 37100 48242 37268 48244
rect 37100 48190 37214 48242
rect 37266 48190 37268 48242
rect 37100 48188 37268 48190
rect 36428 47460 36484 47628
rect 35420 46898 35588 46900
rect 35420 46846 35422 46898
rect 35474 46846 35588 46898
rect 35420 46844 35588 46846
rect 35420 46834 35476 46844
rect 35084 46788 35140 46798
rect 34972 46786 35140 46788
rect 34972 46734 35086 46786
rect 35138 46734 35140 46786
rect 34972 46732 35140 46734
rect 34300 46004 34356 46014
rect 34300 45780 34356 45948
rect 34636 46004 34692 46014
rect 34524 45780 34580 45790
rect 34300 45778 34468 45780
rect 34300 45726 34302 45778
rect 34354 45726 34468 45778
rect 34300 45724 34468 45726
rect 34300 45714 34356 45724
rect 34188 45106 34244 45118
rect 34188 45054 34190 45106
rect 34242 45054 34244 45106
rect 34188 44996 34244 45054
rect 34412 45108 34468 45724
rect 34524 45108 34580 45724
rect 34636 45330 34692 45948
rect 34972 45668 35028 46732
rect 35084 46722 35140 46732
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 46004 35252 46014
rect 35196 45910 35252 45948
rect 35084 45892 35140 45902
rect 35084 45798 35140 45836
rect 34972 45612 35140 45668
rect 34636 45278 34638 45330
rect 34690 45278 34692 45330
rect 34636 45266 34692 45278
rect 34860 45108 34916 45118
rect 34524 45106 34916 45108
rect 34524 45054 34862 45106
rect 34914 45054 34916 45106
rect 34524 45052 34916 45054
rect 34412 45014 34468 45052
rect 34188 44772 34244 44940
rect 33964 44716 34244 44772
rect 33852 43652 33908 43662
rect 33628 43650 33908 43652
rect 33628 43598 33854 43650
rect 33906 43598 33908 43650
rect 33628 43596 33908 43598
rect 33852 43540 33908 43596
rect 33852 43474 33908 43484
rect 33740 42530 33796 42542
rect 33740 42478 33742 42530
rect 33794 42478 33796 42530
rect 33740 42084 33796 42478
rect 33516 42028 33740 42084
rect 33180 41860 33236 41870
rect 33180 41766 33236 41804
rect 33516 41636 33572 42028
rect 33740 41990 33796 42028
rect 33516 41570 33572 41580
rect 33628 41858 33684 41870
rect 33628 41806 33630 41858
rect 33682 41806 33684 41858
rect 33516 41300 33572 41310
rect 33628 41300 33684 41806
rect 33572 41244 33684 41300
rect 33516 41186 33572 41244
rect 33516 41134 33518 41186
rect 33570 41134 33572 41186
rect 33516 41122 33572 41134
rect 33068 41022 33070 41074
rect 33122 41022 33124 41074
rect 33068 41010 33124 41022
rect 33292 40740 33348 40750
rect 33180 40628 33236 40638
rect 32956 39618 33012 39630
rect 32956 39566 32958 39618
rect 33010 39566 33012 39618
rect 32956 39060 33012 39566
rect 33180 39618 33236 40572
rect 33180 39566 33182 39618
rect 33234 39566 33236 39618
rect 33180 39554 33236 39566
rect 33292 40402 33348 40684
rect 33292 40350 33294 40402
rect 33346 40350 33348 40402
rect 32956 38994 33012 39004
rect 33292 39058 33348 40350
rect 33292 39006 33294 39058
rect 33346 39006 33348 39058
rect 33292 38994 33348 39006
rect 33516 40516 33572 40526
rect 33516 38946 33572 40460
rect 33516 38894 33518 38946
rect 33570 38894 33572 38946
rect 33516 38882 33572 38894
rect 33404 38722 33460 38734
rect 33404 38670 33406 38722
rect 33458 38670 33460 38722
rect 33404 38612 33460 38670
rect 33404 38546 33460 38556
rect 32844 38276 32900 38286
rect 33964 38276 34020 44716
rect 34300 44660 34356 44670
rect 34300 43538 34356 44604
rect 34860 44434 34916 45052
rect 34860 44382 34862 44434
rect 34914 44382 34916 44434
rect 34860 44370 34916 44382
rect 34636 44324 34692 44334
rect 34300 43486 34302 43538
rect 34354 43486 34356 43538
rect 34300 43092 34356 43486
rect 34300 43026 34356 43036
rect 34524 44322 34692 44324
rect 34524 44270 34638 44322
rect 34690 44270 34692 44322
rect 34524 44268 34692 44270
rect 34300 42868 34356 42878
rect 34300 42774 34356 42812
rect 34300 42308 34356 42318
rect 34188 42252 34300 42308
rect 34188 42082 34244 42252
rect 34300 42242 34356 42252
rect 34188 42030 34190 42082
rect 34242 42030 34244 42082
rect 34188 42018 34244 42030
rect 34412 42084 34468 42094
rect 34412 41990 34468 42028
rect 34300 41860 34356 41870
rect 34300 41524 34356 41804
rect 34300 41468 34468 41524
rect 34300 41298 34356 41310
rect 34300 41246 34302 41298
rect 34354 41246 34356 41298
rect 34076 41186 34132 41198
rect 34076 41134 34078 41186
rect 34130 41134 34132 41186
rect 34076 40404 34132 41134
rect 34300 40516 34356 41246
rect 34412 41076 34468 41468
rect 34412 40982 34468 41020
rect 34524 40628 34580 44268
rect 34636 44258 34692 44268
rect 34748 43650 34804 43662
rect 34748 43598 34750 43650
rect 34802 43598 34804 43650
rect 34748 43540 34804 43598
rect 34748 43474 34804 43484
rect 34972 43092 35028 43102
rect 34860 42868 34916 42878
rect 34748 42196 34804 42206
rect 34636 42082 34692 42094
rect 34636 42030 34638 42082
rect 34690 42030 34692 42082
rect 34636 41972 34692 42030
rect 34636 41906 34692 41916
rect 34748 41970 34804 42140
rect 34748 41918 34750 41970
rect 34802 41918 34804 41970
rect 34748 41906 34804 41918
rect 34860 41970 34916 42812
rect 34972 42754 35028 43036
rect 34972 42702 34974 42754
rect 35026 42702 35028 42754
rect 34972 42690 35028 42702
rect 35084 42532 35140 45612
rect 35196 44996 35252 45006
rect 35196 44902 35252 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35308 44324 35364 44334
rect 35308 44230 35364 44268
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34860 41918 34862 41970
rect 34914 41918 34916 41970
rect 34300 40422 34356 40460
rect 34412 40572 34580 40628
rect 34076 40338 34132 40348
rect 34188 39844 34244 39854
rect 34188 39750 34244 39788
rect 34412 39058 34468 40572
rect 34860 40292 34916 41918
rect 34860 40226 34916 40236
rect 34972 42476 35140 42532
rect 35196 42866 35252 42878
rect 35196 42814 35198 42866
rect 35250 42814 35252 42866
rect 34412 39006 34414 39058
rect 34466 39006 34468 39058
rect 34412 38994 34468 39006
rect 34636 38834 34692 38846
rect 34636 38782 34638 38834
rect 34690 38782 34692 38834
rect 34636 38668 34692 38782
rect 34972 38668 35028 42476
rect 35196 42194 35252 42814
rect 35196 42142 35198 42194
rect 35250 42142 35252 42194
rect 35196 42130 35252 42142
rect 35308 42420 35364 42430
rect 35308 41972 35364 42364
rect 35308 41748 35364 41916
rect 35532 42196 35588 46844
rect 36204 47404 36484 47460
rect 36540 47460 36596 47470
rect 36204 47346 36260 47404
rect 36540 47366 36596 47404
rect 36204 47294 36206 47346
rect 36258 47294 36260 47346
rect 35868 46116 35924 46126
rect 35868 46022 35924 46060
rect 35756 43650 35812 43662
rect 35756 43598 35758 43650
rect 35810 43598 35812 43650
rect 35644 42644 35700 42654
rect 35644 42550 35700 42588
rect 35756 42420 35812 43598
rect 35868 43538 35924 43550
rect 35868 43486 35870 43538
rect 35922 43486 35924 43538
rect 35868 42868 35924 43486
rect 36204 43426 36260 47294
rect 36316 47236 36372 47246
rect 36316 47142 36372 47180
rect 37100 47236 37156 48188
rect 37212 48178 37268 48188
rect 37212 47460 37268 47470
rect 37212 47366 37268 47404
rect 36988 44324 37044 44334
rect 36988 44230 37044 44268
rect 37100 44100 37156 47180
rect 37324 47068 37380 50428
rect 37660 49924 37716 51100
rect 37884 51156 37940 51166
rect 37884 51062 37940 51100
rect 38332 50708 38388 51324
rect 38556 51380 38612 51998
rect 38780 52052 38836 52062
rect 38780 51490 38836 51996
rect 38780 51438 38782 51490
rect 38834 51438 38836 51490
rect 38780 51426 38836 51438
rect 38556 51314 38612 51324
rect 38332 50642 38388 50652
rect 38780 51156 38836 51166
rect 38780 50594 38836 51100
rect 39004 50708 39060 52108
rect 39116 52098 39172 52108
rect 40572 52162 40628 52174
rect 40572 52110 40574 52162
rect 40626 52110 40628 52162
rect 39452 51940 39508 51950
rect 39900 51940 39956 51950
rect 39452 51846 39508 51884
rect 39564 51938 39956 51940
rect 39564 51886 39902 51938
rect 39954 51886 39956 51938
rect 39564 51884 39956 51886
rect 39452 51604 39508 51614
rect 39564 51604 39620 51884
rect 39900 51874 39956 51884
rect 40124 51938 40180 51950
rect 40124 51886 40126 51938
rect 40178 51886 40180 51938
rect 39452 51602 39620 51604
rect 39452 51550 39454 51602
rect 39506 51550 39620 51602
rect 39452 51548 39620 51550
rect 39452 51538 39508 51548
rect 39004 50642 39060 50652
rect 39116 51380 39172 51390
rect 38780 50542 38782 50594
rect 38834 50542 38836 50594
rect 38780 50530 38836 50542
rect 39004 50484 39060 50494
rect 38892 50372 39060 50428
rect 39116 50428 39172 51324
rect 40012 51380 40068 51390
rect 40124 51380 40180 51886
rect 40068 51324 40180 51380
rect 40572 51380 40628 52110
rect 42028 52162 42084 52174
rect 42028 52110 42030 52162
rect 42082 52110 42084 52162
rect 40796 51940 40852 51950
rect 40796 51846 40852 51884
rect 41020 51940 41076 51950
rect 41020 51938 41188 51940
rect 41020 51886 41022 51938
rect 41074 51886 41188 51938
rect 41020 51884 41188 51886
rect 41020 51874 41076 51884
rect 41020 51716 41076 51726
rect 41020 51602 41076 51660
rect 41020 51550 41022 51602
rect 41074 51550 41076 51602
rect 41020 51538 41076 51550
rect 41132 51490 41188 51884
rect 41132 51438 41134 51490
rect 41186 51438 41188 51490
rect 41132 51380 41188 51438
rect 40572 51324 41076 51380
rect 39228 51156 39284 51166
rect 39228 50706 39284 51100
rect 39228 50654 39230 50706
rect 39282 50654 39284 50706
rect 39228 50642 39284 50654
rect 39788 50708 39844 50718
rect 39340 50596 39396 50606
rect 39340 50502 39396 50540
rect 39116 50372 39396 50428
rect 38108 50036 38164 50046
rect 38108 49942 38164 49980
rect 37660 49858 37716 49868
rect 37436 49810 37492 49822
rect 37436 49758 37438 49810
rect 37490 49758 37492 49810
rect 37436 49700 37492 49758
rect 37436 49634 37492 49644
rect 37884 49810 37940 49822
rect 37884 49758 37886 49810
rect 37938 49758 37940 49810
rect 37884 49028 37940 49758
rect 37996 49700 38052 49710
rect 37996 49606 38052 49644
rect 37884 48962 37940 48972
rect 38444 49028 38500 49038
rect 37772 48804 37828 48814
rect 37772 48802 38052 48804
rect 37772 48750 37774 48802
rect 37826 48750 38052 48802
rect 37772 48748 38052 48750
rect 37772 48738 37828 48748
rect 37996 48354 38052 48748
rect 38444 48466 38500 48972
rect 38444 48414 38446 48466
rect 38498 48414 38500 48466
rect 38444 48402 38500 48414
rect 38892 48468 38948 50372
rect 39004 49140 39060 49150
rect 39004 48804 39060 49084
rect 39004 48738 39060 48748
rect 38892 48412 39060 48468
rect 37996 48302 37998 48354
rect 38050 48302 38052 48354
rect 37436 47684 37492 47694
rect 37436 47570 37492 47628
rect 37436 47518 37438 47570
rect 37490 47518 37492 47570
rect 37436 47506 37492 47518
rect 37660 47572 37716 47582
rect 37324 47012 37492 47068
rect 37324 44548 37380 44558
rect 37324 44454 37380 44492
rect 36988 44044 37156 44100
rect 37324 44324 37380 44334
rect 37436 44324 37492 47012
rect 37324 44322 37492 44324
rect 37324 44270 37326 44322
rect 37378 44270 37492 44322
rect 37324 44268 37492 44270
rect 36204 43374 36206 43426
rect 36258 43374 36260 43426
rect 36204 43362 36260 43374
rect 36316 43540 36372 43550
rect 35868 42802 35924 42812
rect 36316 42754 36372 43484
rect 36316 42702 36318 42754
rect 36370 42702 36372 42754
rect 36316 42690 36372 42702
rect 35756 42354 35812 42364
rect 35980 42642 36036 42654
rect 35980 42590 35982 42642
rect 36034 42590 36036 42642
rect 35868 42196 35924 42206
rect 35532 42194 35924 42196
rect 35532 42142 35870 42194
rect 35922 42142 35924 42194
rect 35532 42140 35924 42142
rect 35532 41970 35588 42140
rect 35868 42130 35924 42140
rect 35980 42196 36036 42590
rect 36092 42532 36148 42542
rect 36092 42530 36372 42532
rect 36092 42478 36094 42530
rect 36146 42478 36372 42530
rect 36092 42476 36372 42478
rect 36092 42466 36148 42476
rect 35980 42130 36036 42140
rect 35532 41918 35534 41970
rect 35586 41918 35588 41970
rect 35532 41906 35588 41918
rect 36204 41970 36260 41982
rect 36204 41918 36206 41970
rect 36258 41918 36260 41970
rect 35308 41692 35588 41748
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35084 41076 35140 41086
rect 35084 40982 35140 41020
rect 35532 41076 35588 41692
rect 36204 41412 36260 41918
rect 35868 41410 36260 41412
rect 35868 41358 36206 41410
rect 36258 41358 36260 41410
rect 35868 41356 36260 41358
rect 35756 41298 35812 41310
rect 35756 41246 35758 41298
rect 35810 41246 35812 41298
rect 35532 41074 35700 41076
rect 35532 41022 35534 41074
rect 35586 41022 35700 41074
rect 35532 41020 35700 41022
rect 35532 41010 35588 41020
rect 35644 40626 35700 41020
rect 35644 40574 35646 40626
rect 35698 40574 35700 40626
rect 35644 40562 35700 40574
rect 35756 40628 35812 41246
rect 35868 41186 35924 41356
rect 36204 41346 36260 41356
rect 35868 41134 35870 41186
rect 35922 41134 35924 41186
rect 35868 41122 35924 41134
rect 36316 41074 36372 42476
rect 36316 41022 36318 41074
rect 36370 41022 36372 41074
rect 36316 40740 36372 41022
rect 36316 40684 36708 40740
rect 35756 40572 36596 40628
rect 35084 40290 35140 40302
rect 35084 40238 35086 40290
rect 35138 40238 35140 40290
rect 35084 39844 35140 40238
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39778 35140 39788
rect 35980 39618 36036 40572
rect 36540 40514 36596 40572
rect 36540 40462 36542 40514
rect 36594 40462 36596 40514
rect 36540 40450 36596 40462
rect 35980 39566 35982 39618
rect 36034 39566 36036 39618
rect 35980 39554 36036 39566
rect 36316 40292 36372 40302
rect 36316 39618 36372 40236
rect 36316 39566 36318 39618
rect 36370 39566 36372 39618
rect 36316 39554 36372 39566
rect 36428 39508 36484 39518
rect 36428 39414 36484 39452
rect 34300 38610 34356 38622
rect 34636 38612 34804 38668
rect 34300 38558 34302 38610
rect 34354 38558 34356 38610
rect 33964 38220 34132 38276
rect 32844 38050 32900 38220
rect 32844 37998 32846 38050
rect 32898 37998 32900 38050
rect 32844 37986 32900 37998
rect 33180 38050 33236 38062
rect 33180 37998 33182 38050
rect 33234 37998 33236 38050
rect 32732 37762 32788 37772
rect 33180 37268 33236 37998
rect 33404 38052 33460 38062
rect 33404 38050 33572 38052
rect 33404 37998 33406 38050
rect 33458 37998 33572 38050
rect 33404 37996 33572 37998
rect 33404 37986 33460 37996
rect 33180 37202 33236 37212
rect 33516 37156 33572 37996
rect 33964 38050 34020 38062
rect 33964 37998 33966 38050
rect 34018 37998 34020 38050
rect 33964 37940 34020 37998
rect 33964 37874 34020 37884
rect 33740 37266 33796 37278
rect 33740 37214 33742 37266
rect 33794 37214 33796 37266
rect 33740 37156 33796 37214
rect 33516 37100 33796 37156
rect 33516 36708 33572 37100
rect 33740 37044 33796 37100
rect 33740 36978 33796 36988
rect 33516 36642 33572 36652
rect 32508 36306 32564 36316
rect 32732 36482 32788 36494
rect 32732 36430 32734 36482
rect 32786 36430 32788 36482
rect 32116 35980 32228 36036
rect 32060 35970 32116 35980
rect 32172 35922 32228 35980
rect 32172 35870 32174 35922
rect 32226 35870 32228 35922
rect 32172 35858 32228 35870
rect 31724 35812 31780 35822
rect 31724 35718 31780 35756
rect 31388 35634 31444 35644
rect 31276 35186 31332 35196
rect 32732 35252 32788 36430
rect 33068 36484 33124 36494
rect 33068 36390 33124 36428
rect 33852 35924 33908 35934
rect 33852 35698 33908 35868
rect 33852 35646 33854 35698
rect 33906 35646 33908 35698
rect 33852 35634 33908 35646
rect 33628 35586 33684 35598
rect 33628 35534 33630 35586
rect 33682 35534 33684 35586
rect 33628 35476 33684 35534
rect 33628 35410 33684 35420
rect 32732 35186 32788 35196
rect 31164 35086 31166 35138
rect 31218 35086 31220 35138
rect 31164 35074 31220 35086
rect 31948 35028 32004 35038
rect 31164 34916 31220 34926
rect 30716 34514 30772 34524
rect 31052 34802 31108 34814
rect 31052 34750 31054 34802
rect 31106 34750 31108 34802
rect 30716 34132 30772 34142
rect 31052 34132 31108 34750
rect 31164 34802 31220 34860
rect 31164 34750 31166 34802
rect 31218 34750 31220 34802
rect 31164 34738 31220 34750
rect 30716 34130 31108 34132
rect 30716 34078 30718 34130
rect 30770 34078 31108 34130
rect 30716 34076 31108 34078
rect 31164 34580 31220 34590
rect 30716 34020 30772 34076
rect 30716 33954 30772 33964
rect 31164 34018 31220 34524
rect 31164 33966 31166 34018
rect 31218 33966 31220 34018
rect 31164 33954 31220 33966
rect 31836 34242 31892 34254
rect 31836 34190 31838 34242
rect 31890 34190 31892 34242
rect 30940 33348 30996 33358
rect 30380 33346 30772 33348
rect 30380 33294 30382 33346
rect 30434 33294 30772 33346
rect 30380 33292 30772 33294
rect 30380 33282 30436 33292
rect 30716 33234 30772 33292
rect 30940 33254 30996 33292
rect 31500 33348 31556 33358
rect 31836 33348 31892 34190
rect 31500 33346 31892 33348
rect 31500 33294 31502 33346
rect 31554 33294 31892 33346
rect 31500 33292 31892 33294
rect 30716 33182 30718 33234
rect 30770 33182 30772 33234
rect 30716 33170 30772 33182
rect 30380 32788 30436 32798
rect 30380 31948 30436 32732
rect 28028 31714 28084 31724
rect 28588 31892 29540 31948
rect 29596 31892 29988 31948
rect 30268 31892 30436 31948
rect 26460 31554 26740 31556
rect 26460 31502 26462 31554
rect 26514 31502 26740 31554
rect 26460 31500 26740 31502
rect 26460 31444 26516 31500
rect 26124 31388 26516 31444
rect 25788 30996 25844 31006
rect 26124 30996 26180 31388
rect 25788 30994 26180 30996
rect 25788 30942 25790 30994
rect 25842 30942 26180 30994
rect 25788 30940 26180 30942
rect 26572 30994 26628 31006
rect 27020 30996 27076 31006
rect 26572 30942 26574 30994
rect 26626 30942 26628 30994
rect 25788 30930 25844 30940
rect 26236 30884 26292 30894
rect 26236 30882 26404 30884
rect 26236 30830 26238 30882
rect 26290 30830 26404 30882
rect 26236 30828 26404 30830
rect 26236 30818 26292 30828
rect 25340 30604 25732 30660
rect 25340 30434 25396 30604
rect 25340 30382 25342 30434
rect 25394 30382 25396 30434
rect 25340 30370 25396 30382
rect 26348 30436 26404 30828
rect 26460 30436 26516 30446
rect 26348 30434 26516 30436
rect 26348 30382 26462 30434
rect 26514 30382 26516 30434
rect 26348 30380 26516 30382
rect 26460 30370 26516 30380
rect 25116 30258 25172 30268
rect 24556 30046 24558 30098
rect 24610 30046 24612 30098
rect 24556 30034 24612 30046
rect 24668 30044 25004 30100
rect 24444 29988 24500 29998
rect 24444 29894 24500 29932
rect 24668 29650 24724 30044
rect 25004 30034 25060 30044
rect 25452 30212 25508 30222
rect 25116 29988 25172 29998
rect 25116 29894 25172 29932
rect 25228 29986 25284 29998
rect 25228 29934 25230 29986
rect 25282 29934 25284 29986
rect 24668 29598 24670 29650
rect 24722 29598 24724 29650
rect 24668 29586 24724 29598
rect 24332 29138 24388 29148
rect 24668 29092 24724 29102
rect 24220 28924 24500 28980
rect 23772 28690 23828 28700
rect 24444 28754 24500 28924
rect 24444 28702 24446 28754
rect 24498 28702 24500 28754
rect 24444 28690 24500 28702
rect 23548 28478 23550 28530
rect 23602 28478 23604 28530
rect 23548 28466 23604 28478
rect 23212 28366 23214 28418
rect 23266 28366 23268 28418
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 28018 19684 28028
rect 23212 28082 23268 28366
rect 23212 28030 23214 28082
rect 23266 28030 23268 28082
rect 23212 28018 23268 28030
rect 24668 28084 24724 29036
rect 25004 28644 25060 28654
rect 25228 28644 25284 29934
rect 25452 29650 25508 30156
rect 25788 30100 25844 30110
rect 25788 30006 25844 30044
rect 25452 29598 25454 29650
rect 25506 29598 25508 29650
rect 25452 29586 25508 29598
rect 25900 28756 25956 28766
rect 25340 28644 25396 28654
rect 25228 28642 25396 28644
rect 25228 28590 25342 28642
rect 25394 28590 25396 28642
rect 25228 28588 25396 28590
rect 25004 28550 25060 28588
rect 25340 28578 25396 28588
rect 25564 28644 25620 28654
rect 24668 27990 24724 28028
rect 25564 28082 25620 28588
rect 25564 28030 25566 28082
rect 25618 28030 25620 28082
rect 25564 28018 25620 28030
rect 25676 28420 25732 28430
rect 19404 27972 19460 27982
rect 19404 27858 19460 27916
rect 22876 27972 22932 27982
rect 22876 27970 23156 27972
rect 22876 27918 22878 27970
rect 22930 27918 23156 27970
rect 22876 27916 23156 27918
rect 22876 27906 22932 27916
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19404 27794 19460 27806
rect 21756 27748 21812 27758
rect 18956 26852 19124 26908
rect 19180 27634 19236 27646
rect 19180 27582 19182 27634
rect 19234 27582 19236 27634
rect 18172 25442 18228 25452
rect 18284 25506 18340 25518
rect 18284 25454 18286 25506
rect 18338 25454 18340 25506
rect 16044 25396 16100 25406
rect 16044 25302 16100 25340
rect 16604 25394 16660 25406
rect 16604 25342 16606 25394
rect 16658 25342 16660 25394
rect 16604 25284 16660 25342
rect 16604 25218 16660 25228
rect 17612 25282 17668 25294
rect 17612 25230 17614 25282
rect 17666 25230 17668 25282
rect 15484 24882 15540 24892
rect 16380 24724 16436 24734
rect 15932 24722 16436 24724
rect 15932 24670 16382 24722
rect 16434 24670 16436 24722
rect 15932 24668 16436 24670
rect 15932 24050 15988 24668
rect 15932 23998 15934 24050
rect 15986 23998 15988 24050
rect 15932 23986 15988 23998
rect 16268 24498 16324 24510
rect 16268 24446 16270 24498
rect 16322 24446 16324 24498
rect 16268 24050 16324 24446
rect 16268 23998 16270 24050
rect 16322 23998 16324 24050
rect 15372 23886 15374 23938
rect 15426 23886 15428 23938
rect 15372 23874 15428 23886
rect 15036 23714 15092 23726
rect 15036 23662 15038 23714
rect 15090 23662 15092 23714
rect 15036 23380 15092 23662
rect 16268 23492 16324 23998
rect 16268 23426 16324 23436
rect 14812 23324 14980 23380
rect 15036 23324 15428 23380
rect 14588 22990 14590 23042
rect 14642 22990 14644 23042
rect 14588 22978 14644 22990
rect 14588 22372 14644 22382
rect 14588 22278 14644 22316
rect 14476 21476 14532 21486
rect 14476 20690 14532 21420
rect 14700 21476 14756 21486
rect 14700 21382 14756 21420
rect 14476 20638 14478 20690
rect 14530 20638 14532 20690
rect 14476 20242 14532 20638
rect 14476 20190 14478 20242
rect 14530 20190 14532 20242
rect 14476 20178 14532 20190
rect 14812 20356 14868 20366
rect 14588 20018 14644 20030
rect 14588 19966 14590 20018
rect 14642 19966 14644 20018
rect 14588 19908 14644 19966
rect 14476 19796 14532 19806
rect 14364 19740 14476 19796
rect 14476 18562 14532 19740
rect 14476 18510 14478 18562
rect 14530 18510 14532 18562
rect 13916 17614 13918 17666
rect 13970 17614 13972 17666
rect 13916 17444 13972 17614
rect 14364 17666 14420 17678
rect 14364 17614 14366 17666
rect 14418 17614 14420 17666
rect 14364 17556 14420 17614
rect 14364 17490 14420 17500
rect 13916 17378 13972 17388
rect 13804 16930 13860 16940
rect 14028 16884 14084 16894
rect 13916 16882 14084 16884
rect 13916 16830 14030 16882
rect 14082 16830 14084 16882
rect 13916 16828 14084 16830
rect 14476 16884 14532 18510
rect 14588 18004 14644 19852
rect 14812 19458 14868 20300
rect 14924 19796 14980 23324
rect 15372 22484 15428 23324
rect 16268 23156 16324 23166
rect 16268 23062 16324 23100
rect 15372 22370 15428 22428
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 15372 22306 15428 22318
rect 16044 22482 16100 22494
rect 16044 22430 16046 22482
rect 16098 22430 16100 22482
rect 15148 22260 15204 22270
rect 15148 22166 15204 22204
rect 15820 22260 15876 22270
rect 15484 21700 15540 21710
rect 15148 21588 15204 21598
rect 15148 21494 15204 21532
rect 15484 20244 15540 21644
rect 15484 20018 15540 20188
rect 15484 19966 15486 20018
rect 15538 19966 15540 20018
rect 15484 19954 15540 19966
rect 15596 21474 15652 21486
rect 15596 21422 15598 21474
rect 15650 21422 15652 21474
rect 15148 19796 15204 19806
rect 14924 19794 15316 19796
rect 14924 19742 15150 19794
rect 15202 19742 15316 19794
rect 14924 19740 15316 19742
rect 15148 19702 15204 19740
rect 14812 19406 14814 19458
rect 14866 19406 14868 19458
rect 14812 19394 14868 19406
rect 15148 19460 15204 19470
rect 14812 18452 14868 18462
rect 14812 18358 14868 18396
rect 14588 17938 14644 17948
rect 14700 18226 14756 18238
rect 14700 18174 14702 18226
rect 14754 18174 14756 18226
rect 14700 17780 14756 18174
rect 14588 16884 14644 16894
rect 14476 16828 14588 16884
rect 13804 16772 13860 16782
rect 13804 16678 13860 16716
rect 13916 16324 13972 16828
rect 14028 16818 14084 16828
rect 14588 16818 14644 16828
rect 14140 16772 14196 16782
rect 14140 16548 14196 16716
rect 14140 16482 14196 16492
rect 14700 16324 14756 17724
rect 13692 15586 13748 15596
rect 13804 16268 13972 16324
rect 14252 16268 14756 16324
rect 15036 17108 15092 17118
rect 13580 15092 13748 15148
rect 13468 14644 13524 14654
rect 13468 14530 13524 14588
rect 13468 14478 13470 14530
rect 13522 14478 13524 14530
rect 13468 14466 13524 14478
rect 13692 14420 13748 15092
rect 13804 15092 13860 16268
rect 14140 16212 14196 16222
rect 13804 15026 13860 15036
rect 13916 16210 14196 16212
rect 13916 16158 14142 16210
rect 14194 16158 14196 16210
rect 13916 16156 14196 16158
rect 13244 12178 13412 12180
rect 13244 12126 13246 12178
rect 13298 12126 13412 12178
rect 13244 12124 13412 12126
rect 13580 12516 13636 12526
rect 13580 12178 13636 12460
rect 13692 12290 13748 14364
rect 13804 14308 13860 14318
rect 13804 13074 13860 14252
rect 13804 13022 13806 13074
rect 13858 13022 13860 13074
rect 13804 13010 13860 13022
rect 13692 12238 13694 12290
rect 13746 12238 13748 12290
rect 13692 12226 13748 12238
rect 13580 12126 13582 12178
rect 13634 12126 13636 12178
rect 13244 10612 13300 12124
rect 13580 12114 13636 12126
rect 13692 11620 13748 11630
rect 13692 11394 13748 11564
rect 13692 11342 13694 11394
rect 13746 11342 13748 11394
rect 13692 11330 13748 11342
rect 13244 10546 13300 10556
rect 13804 10948 13860 10958
rect 13356 10164 13412 10174
rect 13132 10108 13300 10164
rect 13132 9604 13188 9614
rect 13132 9042 13188 9548
rect 13132 8990 13134 9042
rect 13186 8990 13188 9042
rect 13132 8978 13188 8990
rect 12964 8428 13076 8484
rect 12908 8418 12964 8428
rect 12796 8370 12852 8382
rect 12796 8318 12798 8370
rect 12850 8318 12852 8370
rect 12796 8148 12852 8318
rect 12796 8082 12852 8092
rect 13020 8258 13076 8270
rect 13020 8206 13022 8258
rect 13074 8206 13076 8258
rect 12684 7534 12686 7586
rect 12738 7534 12740 7586
rect 12684 6580 12740 7534
rect 13020 7476 13076 8206
rect 13244 7700 13300 10108
rect 13412 10108 13524 10164
rect 13356 10098 13412 10108
rect 13356 8932 13412 8942
rect 13356 8838 13412 8876
rect 13356 8260 13412 8270
rect 13468 8260 13524 10108
rect 13692 10050 13748 10062
rect 13692 9998 13694 10050
rect 13746 9998 13748 10050
rect 13692 9940 13748 9998
rect 13692 9874 13748 9884
rect 13804 9826 13860 10892
rect 13916 10834 13972 16156
rect 14140 16146 14196 16156
rect 14252 15876 14308 16268
rect 14588 16100 14644 16110
rect 14812 16100 14868 16110
rect 14588 16098 14812 16100
rect 14588 16046 14590 16098
rect 14642 16046 14812 16098
rect 14588 16044 14812 16046
rect 14588 16034 14644 16044
rect 14812 16034 14868 16044
rect 14140 15820 14308 15876
rect 14924 15986 14980 15998
rect 14924 15934 14926 15986
rect 14978 15934 14980 15986
rect 14028 13748 14084 13758
rect 14028 13186 14084 13692
rect 14028 13134 14030 13186
rect 14082 13134 14084 13186
rect 14028 13122 14084 13134
rect 14028 12066 14084 12078
rect 14028 12014 14030 12066
rect 14082 12014 14084 12066
rect 14028 11844 14084 12014
rect 14028 11778 14084 11788
rect 13916 10782 13918 10834
rect 13970 10782 13972 10834
rect 13916 10770 13972 10782
rect 14028 11506 14084 11518
rect 14028 11454 14030 11506
rect 14082 11454 14084 11506
rect 14028 11060 14084 11454
rect 14028 10724 14084 11004
rect 14028 10658 14084 10668
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13804 9762 13860 9774
rect 13916 10388 13972 10398
rect 13580 9716 13636 9726
rect 13580 8708 13636 9660
rect 13692 9602 13748 9614
rect 13692 9550 13694 9602
rect 13746 9550 13748 9602
rect 13692 9380 13748 9550
rect 13692 9314 13748 9324
rect 13692 9154 13748 9166
rect 13692 9102 13694 9154
rect 13746 9102 13748 9154
rect 13692 9044 13748 9102
rect 13692 8978 13748 8988
rect 13580 8652 13748 8708
rect 13356 8258 13524 8260
rect 13356 8206 13358 8258
rect 13410 8206 13524 8258
rect 13356 8204 13524 8206
rect 13580 8484 13636 8494
rect 13580 8260 13636 8428
rect 13356 8194 13412 8204
rect 13580 8146 13636 8204
rect 13692 8258 13748 8652
rect 13692 8206 13694 8258
rect 13746 8206 13748 8258
rect 13692 8194 13748 8206
rect 13580 8094 13582 8146
rect 13634 8094 13636 8146
rect 13580 8082 13636 8094
rect 13804 8036 13860 8046
rect 12236 6130 12404 6132
rect 12236 6078 12238 6130
rect 12290 6078 12404 6130
rect 12236 6076 12404 6078
rect 12572 6132 12628 6142
rect 12236 6066 12292 6076
rect 11228 4562 11508 4564
rect 11228 4510 11230 4562
rect 11282 4510 11508 4562
rect 11228 4508 11508 4510
rect 11564 5236 11620 5246
rect 11228 4498 11284 4508
rect 10892 3614 10894 3666
rect 10946 3614 10948 3666
rect 10892 3602 10948 3614
rect 11564 3668 11620 5180
rect 11788 5012 11844 5022
rect 11564 3602 11620 3612
rect 11676 4226 11732 4238
rect 11676 4174 11678 4226
rect 11730 4174 11732 4226
rect 10780 3266 10836 3276
rect 11340 3330 11396 3342
rect 11340 3278 11342 3330
rect 11394 3278 11396 3330
rect 8988 3154 9044 3164
rect 8316 2818 8372 2828
rect 11340 2548 11396 3278
rect 11676 3108 11732 4174
rect 11788 3666 11844 4956
rect 11900 4452 11956 4462
rect 11900 4358 11956 4396
rect 11788 3614 11790 3666
rect 11842 3614 11844 3666
rect 11788 3602 11844 3614
rect 12124 3668 12180 5852
rect 12572 5906 12628 6076
rect 12572 5854 12574 5906
rect 12626 5854 12628 5906
rect 12572 5842 12628 5854
rect 12684 5348 12740 6524
rect 12796 7420 13020 7476
rect 12796 6130 12852 7420
rect 13020 7410 13076 7420
rect 13132 7588 13188 7598
rect 12908 6916 12964 6926
rect 12908 6690 12964 6860
rect 12908 6638 12910 6690
rect 12962 6638 12964 6690
rect 12908 6468 12964 6638
rect 13132 6580 13188 7532
rect 13244 6804 13300 7644
rect 13244 6738 13300 6748
rect 13356 7812 13412 7822
rect 13356 7474 13412 7756
rect 13804 7586 13860 7980
rect 13804 7534 13806 7586
rect 13858 7534 13860 7586
rect 13804 7522 13860 7534
rect 13916 7588 13972 10332
rect 14140 10164 14196 15820
rect 14812 15652 14868 15662
rect 14588 15540 14644 15550
rect 14476 15202 14532 15214
rect 14476 15150 14478 15202
rect 14530 15150 14532 15202
rect 14476 15092 14532 15150
rect 14476 15026 14532 15036
rect 14588 14642 14644 15484
rect 14588 14590 14590 14642
rect 14642 14590 14644 14642
rect 14476 14308 14532 14318
rect 14476 13858 14532 14252
rect 14588 13972 14644 14590
rect 14588 13906 14644 13916
rect 14700 15090 14756 15102
rect 14700 15038 14702 15090
rect 14754 15038 14756 15090
rect 14476 13806 14478 13858
rect 14530 13806 14532 13858
rect 14476 13794 14532 13806
rect 14700 13748 14756 15038
rect 14700 13654 14756 13692
rect 14252 13076 14308 13086
rect 14252 10276 14308 13020
rect 14476 13076 14532 13086
rect 14364 12964 14420 12974
rect 14364 12870 14420 12908
rect 14252 10210 14308 10220
rect 14476 10834 14532 13020
rect 14588 12740 14644 12750
rect 14588 12178 14644 12684
rect 14812 12404 14868 15596
rect 14924 14532 14980 15934
rect 15036 15988 15092 17052
rect 15148 16100 15204 19404
rect 15260 18562 15316 19740
rect 15596 19460 15652 21422
rect 15820 20802 15876 22204
rect 16044 22036 16100 22430
rect 16380 22372 16436 24668
rect 17388 24724 17444 24734
rect 16492 23940 16548 23950
rect 16492 23846 16548 23884
rect 16492 23604 16548 23614
rect 16492 22594 16548 23548
rect 17388 23378 17444 24668
rect 17612 24388 17668 25230
rect 18284 25172 18340 25454
rect 18732 25508 18788 25518
rect 18732 25414 18788 25452
rect 18172 25116 18340 25172
rect 17836 24948 17892 24958
rect 17836 24722 17892 24892
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24658 17892 24670
rect 17612 24322 17668 24332
rect 18060 24388 18116 24398
rect 17388 23326 17390 23378
rect 17442 23326 17444 23378
rect 17388 23314 17444 23326
rect 16716 23268 16772 23278
rect 16716 23154 16772 23212
rect 16716 23102 16718 23154
rect 16770 23102 16772 23154
rect 16716 23090 16772 23102
rect 17948 23044 18004 23054
rect 16492 22542 16494 22594
rect 16546 22542 16548 22594
rect 16492 22530 16548 22542
rect 17724 23042 18004 23044
rect 17724 22990 17950 23042
rect 18002 22990 18004 23042
rect 17724 22988 18004 22990
rect 16044 21970 16100 21980
rect 16156 22316 16380 22372
rect 16044 21812 16100 21822
rect 16156 21812 16212 22316
rect 16380 22278 16436 22316
rect 17164 22484 17220 22494
rect 17164 22370 17220 22428
rect 17164 22318 17166 22370
rect 17218 22318 17220 22370
rect 16716 21924 16772 21934
rect 16044 21810 16212 21812
rect 16044 21758 16046 21810
rect 16098 21758 16212 21810
rect 16044 21756 16212 21758
rect 16492 21812 16548 21822
rect 16044 21746 16100 21756
rect 15820 20750 15822 20802
rect 15874 20750 15876 20802
rect 15820 20738 15876 20750
rect 16044 21588 16100 21598
rect 15932 20690 15988 20702
rect 15932 20638 15934 20690
rect 15986 20638 15988 20690
rect 15596 19394 15652 19404
rect 15708 20244 15764 20254
rect 15708 20018 15764 20188
rect 15708 19966 15710 20018
rect 15762 19966 15764 20018
rect 15260 18510 15262 18562
rect 15314 18510 15316 18562
rect 15260 17668 15316 18510
rect 15260 17602 15316 17612
rect 15484 19236 15540 19246
rect 15708 19236 15764 19966
rect 15484 19234 15764 19236
rect 15484 19182 15486 19234
rect 15538 19182 15764 19234
rect 15484 19180 15764 19182
rect 15484 17444 15540 19180
rect 15148 16034 15204 16044
rect 15260 17388 15540 17444
rect 15708 18004 15764 18014
rect 15036 15922 15092 15932
rect 15036 15428 15092 15438
rect 15036 15202 15092 15372
rect 15260 15314 15316 17388
rect 15484 16884 15540 16894
rect 15372 16212 15428 16222
rect 15372 16098 15428 16156
rect 15372 16046 15374 16098
rect 15426 16046 15428 16098
rect 15372 16034 15428 16046
rect 15260 15262 15262 15314
rect 15314 15262 15316 15314
rect 15260 15250 15316 15262
rect 15372 15652 15428 15662
rect 15036 15150 15038 15202
rect 15090 15150 15092 15202
rect 15036 15138 15092 15150
rect 15372 15148 15428 15596
rect 14924 14466 14980 14476
rect 15260 15092 15428 15148
rect 15484 15148 15540 16828
rect 15708 16882 15764 17948
rect 15820 17668 15876 17678
rect 15820 17332 15876 17612
rect 15820 17266 15876 17276
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16818 15764 16830
rect 15596 16548 15652 16558
rect 15596 15540 15652 16492
rect 15820 16100 15876 16110
rect 15596 15474 15652 15484
rect 15708 16044 15820 16100
rect 15484 15092 15652 15148
rect 14924 13524 14980 13534
rect 14924 12740 14980 13468
rect 15260 13524 15316 15092
rect 15372 14644 15428 14654
rect 15372 14084 15428 14588
rect 15372 14018 15428 14028
rect 15260 13458 15316 13468
rect 15484 13970 15540 13982
rect 15484 13918 15486 13970
rect 15538 13918 15540 13970
rect 15484 13524 15540 13918
rect 15596 13972 15652 15092
rect 15596 13906 15652 13916
rect 15484 13458 15540 13468
rect 15596 13746 15652 13758
rect 15596 13694 15598 13746
rect 15650 13694 15652 13746
rect 15036 12964 15092 12974
rect 15036 12870 15092 12908
rect 14924 12684 15092 12740
rect 14812 12348 14980 12404
rect 14812 12180 14868 12190
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 14588 12114 14644 12126
rect 14700 12178 14868 12180
rect 14700 12126 14814 12178
rect 14866 12126 14868 12178
rect 14700 12124 14868 12126
rect 14476 10782 14478 10834
rect 14530 10782 14532 10834
rect 14140 10098 14196 10108
rect 14364 10052 14420 10062
rect 14364 9826 14420 9996
rect 14364 9774 14366 9826
rect 14418 9774 14420 9826
rect 14364 9716 14420 9774
rect 14476 9828 14532 10782
rect 14588 11732 14644 11742
rect 14588 10388 14644 11676
rect 14588 10322 14644 10332
rect 14700 11284 14756 12124
rect 14812 12114 14868 12124
rect 14700 9938 14756 11228
rect 14812 11954 14868 11966
rect 14812 11902 14814 11954
rect 14866 11902 14868 11954
rect 14812 10948 14868 11902
rect 14924 11732 14980 12348
rect 14924 11666 14980 11676
rect 14812 10882 14868 10892
rect 14924 11394 14980 11406
rect 14924 11342 14926 11394
rect 14978 11342 14980 11394
rect 14924 10612 14980 11342
rect 15036 11060 15092 12684
rect 15596 12292 15652 13694
rect 15596 12226 15652 12236
rect 15036 10994 15092 11004
rect 14924 10546 14980 10556
rect 15260 10610 15316 10622
rect 15260 10558 15262 10610
rect 15314 10558 15316 10610
rect 15036 10500 15092 10510
rect 15036 10498 15204 10500
rect 15036 10446 15038 10498
rect 15090 10446 15204 10498
rect 15036 10444 15204 10446
rect 15036 10434 15092 10444
rect 14924 10276 14980 10286
rect 14700 9886 14702 9938
rect 14754 9886 14756 9938
rect 14700 9874 14756 9886
rect 14812 10164 14868 10174
rect 14476 9762 14532 9772
rect 13916 7522 13972 7532
rect 14028 9660 14420 9716
rect 14588 9716 14644 9726
rect 13356 7422 13358 7474
rect 13410 7422 13412 7474
rect 13356 6580 13412 7422
rect 13468 7476 13524 7486
rect 13468 7382 13524 7420
rect 13692 7252 13748 7262
rect 13692 6916 13748 7196
rect 13132 6524 13300 6580
rect 12908 6402 12964 6412
rect 12796 6078 12798 6130
rect 12850 6078 12852 6130
rect 12796 6066 12852 6078
rect 12684 5282 12740 5292
rect 13244 5906 13300 6524
rect 13356 6514 13412 6524
rect 13468 6860 13748 6916
rect 14028 6914 14084 9660
rect 14140 9156 14196 9194
rect 14140 9090 14196 9100
rect 14588 9042 14644 9660
rect 14588 8990 14590 9042
rect 14642 8990 14644 9042
rect 14588 8978 14644 8990
rect 14476 8372 14532 8382
rect 14700 8372 14756 8382
rect 14532 8316 14644 8372
rect 14476 8306 14532 8316
rect 14588 8258 14644 8316
rect 14700 8278 14756 8316
rect 14588 8206 14590 8258
rect 14642 8206 14644 8258
rect 14588 8194 14644 8206
rect 14812 8260 14868 10108
rect 14924 9266 14980 10220
rect 15148 9492 15204 10444
rect 15260 10388 15316 10558
rect 15596 10610 15652 10622
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15260 10322 15316 10332
rect 15484 10498 15540 10510
rect 15484 10446 15486 10498
rect 15538 10446 15540 10498
rect 15372 10052 15428 10062
rect 15372 9828 15428 9996
rect 15372 9762 15428 9772
rect 15484 9716 15540 10446
rect 15484 9650 15540 9660
rect 15260 9492 15316 9502
rect 15148 9436 15260 9492
rect 15260 9426 15316 9436
rect 14924 9214 14926 9266
rect 14978 9214 14980 9266
rect 14924 9202 14980 9214
rect 14924 9044 14980 9054
rect 15596 9044 15652 10558
rect 14924 8950 14980 8988
rect 15260 8988 15652 9044
rect 15260 8428 15316 8988
rect 15484 8820 15540 8830
rect 15036 8372 15316 8428
rect 15372 8596 15428 8606
rect 14924 8260 14980 8270
rect 14812 8258 14980 8260
rect 14812 8206 14926 8258
rect 14978 8206 14980 8258
rect 14812 8204 14980 8206
rect 14140 8148 14196 8158
rect 14476 8148 14532 8158
rect 14196 8146 14532 8148
rect 14196 8094 14478 8146
rect 14530 8094 14532 8146
rect 14196 8092 14532 8094
rect 14140 8082 14196 8092
rect 14476 7924 14532 8092
rect 14476 7868 14756 7924
rect 14028 6862 14030 6914
rect 14082 6862 14084 6914
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 13244 5236 13300 5854
rect 13468 5572 13524 6860
rect 14028 6850 14084 6862
rect 14140 7474 14196 7486
rect 14140 7422 14142 7474
rect 14194 7422 14196 7474
rect 13244 5170 13300 5180
rect 13356 5516 13524 5572
rect 13580 6690 13636 6702
rect 13580 6638 13582 6690
rect 13634 6638 13636 6690
rect 12236 5124 12292 5134
rect 13356 5124 13412 5516
rect 13468 5348 13524 5358
rect 13468 5254 13524 5292
rect 13580 5124 13636 6638
rect 14028 6692 14084 6702
rect 14028 6598 14084 6636
rect 13692 6580 13748 6590
rect 13692 5906 13748 6524
rect 13692 5854 13694 5906
rect 13746 5854 13748 5906
rect 13692 5796 13748 5854
rect 13692 5730 13748 5740
rect 13916 5906 13972 5918
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 13804 5684 13860 5694
rect 13692 5236 13748 5246
rect 13692 5142 13748 5180
rect 13356 5068 13524 5124
rect 12236 5030 12292 5068
rect 12572 4900 12628 4910
rect 12572 4806 12628 4844
rect 13356 4788 13412 4798
rect 12684 4676 12740 4686
rect 12236 4450 12292 4462
rect 12236 4398 12238 4450
rect 12290 4398 12292 4450
rect 12236 4340 12292 4398
rect 12236 4274 12292 4284
rect 12684 3778 12740 4620
rect 12908 4340 12964 4350
rect 12908 4246 12964 4284
rect 13356 4338 13412 4732
rect 13356 4286 13358 4338
rect 13410 4286 13412 4338
rect 13356 4274 13412 4286
rect 12684 3726 12686 3778
rect 12738 3726 12740 3778
rect 12236 3668 12292 3678
rect 12124 3666 12292 3668
rect 12124 3614 12238 3666
rect 12290 3614 12292 3666
rect 12124 3612 12292 3614
rect 12236 3602 12292 3612
rect 12684 3666 12740 3726
rect 12684 3614 12686 3666
rect 12738 3614 12740 3666
rect 12684 3602 12740 3614
rect 13356 3892 13412 3902
rect 13356 3666 13412 3836
rect 13356 3614 13358 3666
rect 13410 3614 13412 3666
rect 13356 3602 13412 3614
rect 13468 3556 13524 5068
rect 13580 5058 13636 5068
rect 13692 4564 13748 4574
rect 13692 4470 13748 4508
rect 13804 3666 13860 5628
rect 13916 5572 13972 5854
rect 14140 5794 14196 7422
rect 14700 7362 14756 7868
rect 14700 7310 14702 7362
rect 14754 7310 14756 7362
rect 14700 7298 14756 7310
rect 14476 6018 14532 6030
rect 14476 5966 14478 6018
rect 14530 5966 14532 6018
rect 14140 5742 14142 5794
rect 14194 5742 14196 5794
rect 14140 5730 14196 5742
rect 14252 5906 14308 5918
rect 14252 5854 14254 5906
rect 14306 5854 14308 5906
rect 13916 5506 13972 5516
rect 14252 5348 14308 5854
rect 14476 5796 14532 5966
rect 14476 5730 14532 5740
rect 14700 5906 14756 5918
rect 14700 5854 14702 5906
rect 14754 5854 14756 5906
rect 13916 5292 14252 5348
rect 13916 4898 13972 5292
rect 14252 5254 14308 5292
rect 14476 5236 14532 5246
rect 14028 5124 14084 5134
rect 14476 5124 14532 5180
rect 14028 5122 14532 5124
rect 14028 5070 14030 5122
rect 14082 5070 14532 5122
rect 14028 5068 14532 5070
rect 14028 5058 14084 5068
rect 13916 4846 13918 4898
rect 13970 4846 13972 4898
rect 13916 4788 13972 4846
rect 14140 4900 14196 4910
rect 14140 4806 14196 4844
rect 14700 4788 14756 5854
rect 14812 4900 14868 8204
rect 14924 8194 14980 8204
rect 15036 7476 15092 8372
rect 14924 6692 14980 6702
rect 15036 6692 15092 7420
rect 14924 6690 15092 6692
rect 14924 6638 14926 6690
rect 14978 6638 15092 6690
rect 14924 6636 15092 6638
rect 15148 7474 15204 7486
rect 15148 7422 15150 7474
rect 15202 7422 15204 7474
rect 15148 6916 15204 7422
rect 14924 6626 14980 6636
rect 15036 6020 15092 6030
rect 15036 5906 15092 5964
rect 15036 5854 15038 5906
rect 15090 5854 15092 5906
rect 14924 5236 14980 5246
rect 14924 5122 14980 5180
rect 14924 5070 14926 5122
rect 14978 5070 14980 5122
rect 14924 5058 14980 5070
rect 14812 4898 14980 4900
rect 14812 4846 14814 4898
rect 14866 4846 14980 4898
rect 14812 4844 14980 4846
rect 14812 4834 14868 4844
rect 13916 4722 13972 4732
rect 14252 4732 14756 4788
rect 13804 3614 13806 3666
rect 13858 3614 13860 3666
rect 13804 3602 13860 3614
rect 14140 4452 14196 4462
rect 14140 3668 14196 4396
rect 14252 4338 14308 4732
rect 14252 4286 14254 4338
rect 14306 4286 14308 4338
rect 14252 4274 14308 4286
rect 14700 4116 14756 4732
rect 14812 4340 14868 4350
rect 14812 4246 14868 4284
rect 14700 4050 14756 4060
rect 14140 3574 14196 3612
rect 14252 4004 14308 4014
rect 13468 3490 13524 3500
rect 14252 3444 14308 3948
rect 14252 3378 14308 3388
rect 14588 3444 14644 3482
rect 14588 3378 14644 3388
rect 11676 3042 11732 3052
rect 11340 2482 11396 2492
rect 14924 2772 14980 4844
rect 15036 4004 15092 5854
rect 15148 5572 15204 6860
rect 15260 6468 15316 6478
rect 15260 6374 15316 6412
rect 15372 6244 15428 8540
rect 15484 8148 15540 8764
rect 15708 8260 15764 16044
rect 15820 16006 15876 16044
rect 15820 15876 15876 15886
rect 15820 15538 15876 15820
rect 15820 15486 15822 15538
rect 15874 15486 15876 15538
rect 15820 15204 15876 15486
rect 15820 15138 15876 15148
rect 15932 14756 15988 20638
rect 16044 19122 16100 21532
rect 16492 21586 16548 21756
rect 16492 21534 16494 21586
rect 16546 21534 16548 21586
rect 16268 21364 16324 21374
rect 16044 19070 16046 19122
rect 16098 19070 16100 19122
rect 16044 18452 16100 19070
rect 16044 18358 16100 18396
rect 16156 20020 16212 20030
rect 16156 19124 16212 19964
rect 16156 18564 16212 19068
rect 16156 18228 16212 18508
rect 15820 14700 15988 14756
rect 16044 18172 16212 18228
rect 16268 18228 16324 21308
rect 16492 20244 16548 21534
rect 16492 20178 16548 20188
rect 16380 20018 16436 20030
rect 16380 19966 16382 20018
rect 16434 19966 16436 20018
rect 16380 18564 16436 19966
rect 16604 20020 16660 20030
rect 16604 19926 16660 19964
rect 16380 18498 16436 18508
rect 16268 18172 16436 18228
rect 15820 13074 15876 14700
rect 15932 14532 15988 14570
rect 15932 14466 15988 14476
rect 16044 14196 16100 18172
rect 16268 17444 16324 17454
rect 16268 17350 16324 17388
rect 16156 16770 16212 16782
rect 16156 16718 16158 16770
rect 16210 16718 16212 16770
rect 16156 16660 16212 16718
rect 16156 15876 16212 16604
rect 16156 15810 16212 15820
rect 16268 15764 16324 15774
rect 16268 15428 16324 15708
rect 16268 15334 16324 15372
rect 16380 14532 16436 18172
rect 16492 17220 16548 17230
rect 16492 15092 16548 17164
rect 16716 16212 16772 21868
rect 17164 21812 17220 22318
rect 17276 22372 17332 22382
rect 17276 22258 17332 22316
rect 17276 22206 17278 22258
rect 17330 22206 17332 22258
rect 17276 22194 17332 22206
rect 17500 22146 17556 22158
rect 17500 22094 17502 22146
rect 17554 22094 17556 22146
rect 17500 21924 17556 22094
rect 17500 21858 17556 21868
rect 17388 21812 17444 21822
rect 17164 21810 17444 21812
rect 17164 21758 17390 21810
rect 17442 21758 17444 21810
rect 17164 21756 17444 21758
rect 17388 21746 17444 21756
rect 16828 21698 16884 21710
rect 16828 21646 16830 21698
rect 16882 21646 16884 21698
rect 16828 20916 16884 21646
rect 17388 21252 17444 21262
rect 16828 20860 17332 20916
rect 17164 20692 17220 20702
rect 16828 20132 16884 20142
rect 16828 20038 16884 20076
rect 16940 20020 16996 20030
rect 16940 19926 16996 19964
rect 16940 18676 16996 18686
rect 17164 18676 17220 20636
rect 17276 18788 17332 20860
rect 17388 20802 17444 21196
rect 17388 20750 17390 20802
rect 17442 20750 17444 20802
rect 17388 20356 17444 20750
rect 17724 20804 17780 22988
rect 17948 22978 18004 22988
rect 18060 22484 18116 24332
rect 17948 22428 18116 22484
rect 18172 22484 18228 25116
rect 18284 24948 18340 24958
rect 18732 24948 18788 24958
rect 18340 24892 18452 24948
rect 18284 24882 18340 24892
rect 18396 24388 18452 24892
rect 18788 24892 18900 24948
rect 18732 24882 18788 24892
rect 18508 24610 18564 24622
rect 18508 24558 18510 24610
rect 18562 24558 18564 24610
rect 18508 24500 18564 24558
rect 18732 24500 18788 24510
rect 18508 24498 18788 24500
rect 18508 24446 18734 24498
rect 18786 24446 18788 24498
rect 18508 24444 18788 24446
rect 18396 24332 18564 24388
rect 18284 24164 18340 24174
rect 18284 24070 18340 24108
rect 18508 23378 18564 24332
rect 18620 23940 18676 23950
rect 18620 23604 18676 23884
rect 18620 23538 18676 23548
rect 18732 23380 18788 24444
rect 18508 23326 18510 23378
rect 18562 23326 18564 23378
rect 18508 23314 18564 23326
rect 18620 23324 18788 23380
rect 18172 22428 18452 22484
rect 17948 22260 18004 22428
rect 18172 22260 18228 22270
rect 17948 22258 18228 22260
rect 17948 22206 18174 22258
rect 18226 22206 18228 22258
rect 17948 22204 18228 22206
rect 18060 21700 18116 22204
rect 18172 22194 18228 22204
rect 18284 22260 18340 22270
rect 18284 22166 18340 22204
rect 18060 21634 18116 21644
rect 17948 21588 18004 21598
rect 17948 21494 18004 21532
rect 17724 20748 18340 20804
rect 17388 20290 17444 20300
rect 17836 20580 17892 20590
rect 17724 20020 17780 20030
rect 17724 19926 17780 19964
rect 17836 19572 17892 20524
rect 17612 19516 17892 19572
rect 17500 18788 17556 18798
rect 17276 18732 17500 18788
rect 16940 18562 16996 18620
rect 16940 18510 16942 18562
rect 16994 18510 16996 18562
rect 16940 18498 16996 18510
rect 17052 18620 17220 18676
rect 16716 16146 16772 16156
rect 16828 18004 16884 18014
rect 16828 17666 16884 17948
rect 16828 17614 16830 17666
rect 16882 17614 16884 17666
rect 16716 15540 16772 15550
rect 16604 15316 16660 15326
rect 16604 15222 16660 15260
rect 16492 15026 16548 15036
rect 16716 14642 16772 15484
rect 16828 15426 16884 17614
rect 16828 15374 16830 15426
rect 16882 15374 16884 15426
rect 16828 15362 16884 15374
rect 16716 14590 16718 14642
rect 16770 14590 16772 14642
rect 16716 14578 16772 14590
rect 16380 14476 16660 14532
rect 15820 13022 15822 13074
rect 15874 13022 15876 13074
rect 15820 13010 15876 13022
rect 15932 14140 16100 14196
rect 16268 14418 16324 14430
rect 16268 14366 16270 14418
rect 16322 14366 16324 14418
rect 15932 12178 15988 14140
rect 15932 12126 15934 12178
rect 15986 12126 15988 12178
rect 15932 12114 15988 12126
rect 16044 13972 16100 13982
rect 16044 11788 16100 13916
rect 16268 13634 16324 14366
rect 16268 13582 16270 13634
rect 16322 13582 16324 13634
rect 16268 12964 16324 13582
rect 16268 12898 16324 12908
rect 16268 12292 16324 12302
rect 16268 12198 16324 12236
rect 15820 11732 16100 11788
rect 15820 10610 15876 11732
rect 16268 11396 16324 11406
rect 16268 11394 16436 11396
rect 16268 11342 16270 11394
rect 16322 11342 16436 11394
rect 16268 11340 16436 11342
rect 16268 11330 16324 11340
rect 15820 10558 15822 10610
rect 15874 10558 15876 10610
rect 15820 10500 15876 10558
rect 15820 10434 15876 10444
rect 16268 10498 16324 10510
rect 16268 10446 16270 10498
rect 16322 10446 16324 10498
rect 16268 10164 16324 10446
rect 16268 10098 16324 10108
rect 16156 10052 16212 10062
rect 16156 9958 16212 9996
rect 16044 9826 16100 9838
rect 16044 9774 16046 9826
rect 16098 9774 16100 9826
rect 16044 9604 16100 9774
rect 16044 9538 16100 9548
rect 16156 9492 16212 9502
rect 15932 9044 15988 9054
rect 15932 8950 15988 8988
rect 16156 9044 16212 9436
rect 16156 8930 16212 8988
rect 16156 8878 16158 8930
rect 16210 8878 16212 8930
rect 16156 8866 16212 8878
rect 16268 9042 16324 9054
rect 16268 8990 16270 9042
rect 16322 8990 16324 9042
rect 15708 8204 15988 8260
rect 15484 8092 15652 8148
rect 15484 7586 15540 7598
rect 15484 7534 15486 7586
rect 15538 7534 15540 7586
rect 15484 7476 15540 7534
rect 15484 7410 15540 7420
rect 15596 6914 15652 8092
rect 15932 7700 15988 8204
rect 15820 7698 15988 7700
rect 15820 7646 15934 7698
rect 15986 7646 15988 7698
rect 15820 7644 15988 7646
rect 15708 7588 15764 7598
rect 15708 7494 15764 7532
rect 15596 6862 15598 6914
rect 15650 6862 15652 6914
rect 15596 6850 15652 6862
rect 15820 6692 15876 7644
rect 15932 7634 15988 7644
rect 16044 7924 16100 7934
rect 16044 7474 16100 7868
rect 16044 7422 16046 7474
rect 16098 7422 16100 7474
rect 16044 7252 16100 7422
rect 16044 7186 16100 7196
rect 15372 6178 15428 6188
rect 15484 6636 15876 6692
rect 15932 6802 15988 6814
rect 15932 6750 15934 6802
rect 15986 6750 15988 6802
rect 15932 6692 15988 6750
rect 16156 6692 16212 6702
rect 15932 6690 16212 6692
rect 15932 6638 16158 6690
rect 16210 6638 16212 6690
rect 15932 6636 16212 6638
rect 15148 5506 15204 5516
rect 15260 6018 15316 6030
rect 15260 5966 15262 6018
rect 15314 5966 15316 6018
rect 15148 5236 15204 5246
rect 15148 5142 15204 5180
rect 15260 4452 15316 5966
rect 15372 5682 15428 5694
rect 15372 5630 15374 5682
rect 15426 5630 15428 5682
rect 15372 5122 15428 5630
rect 15372 5070 15374 5122
rect 15426 5070 15428 5122
rect 15372 5058 15428 5070
rect 15260 4386 15316 4396
rect 15260 4228 15316 4238
rect 15484 4228 15540 6636
rect 16156 6626 16212 6636
rect 16268 6580 16324 8990
rect 16380 8372 16436 11340
rect 16492 9268 16548 9278
rect 16492 8932 16548 9212
rect 16492 8866 16548 8876
rect 16380 8306 16436 8316
rect 16492 8260 16548 8270
rect 16380 8146 16436 8158
rect 16380 8094 16382 8146
rect 16434 8094 16436 8146
rect 16380 7476 16436 8094
rect 16380 7410 16436 7420
rect 16492 7140 16548 8204
rect 16492 7074 16548 7084
rect 16604 6916 16660 14476
rect 16828 13748 16884 13758
rect 16716 13692 16828 13748
rect 16716 12178 16772 13692
rect 16828 13654 16884 13692
rect 16716 12126 16718 12178
rect 16770 12126 16772 12178
rect 16716 12114 16772 12126
rect 16940 12964 16996 12974
rect 16828 11844 16884 11854
rect 16716 11732 16772 11742
rect 16716 10610 16772 11676
rect 16828 11394 16884 11788
rect 16828 11342 16830 11394
rect 16882 11342 16884 11394
rect 16828 11330 16884 11342
rect 16940 11508 16996 12908
rect 16716 10558 16718 10610
rect 16770 10558 16772 10610
rect 16716 10546 16772 10558
rect 16828 10500 16884 10510
rect 16716 8820 16772 8830
rect 16716 8726 16772 8764
rect 16828 8148 16884 10444
rect 16828 8082 16884 8092
rect 16940 7700 16996 11452
rect 16828 7644 16940 7700
rect 16828 7586 16884 7644
rect 16940 7634 16996 7644
rect 16828 7534 16830 7586
rect 16882 7534 16884 7586
rect 16828 7522 16884 7534
rect 16828 7364 16884 7374
rect 16268 6514 16324 6524
rect 16380 6860 16660 6916
rect 16716 7308 16828 7364
rect 15820 6466 15876 6478
rect 15820 6414 15822 6466
rect 15874 6414 15876 6466
rect 15596 6020 15652 6030
rect 15596 5122 15652 5964
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 15596 4676 15652 5070
rect 15596 4610 15652 4620
rect 15820 5796 15876 6414
rect 15260 4226 15484 4228
rect 15260 4174 15262 4226
rect 15314 4174 15484 4226
rect 15260 4172 15484 4174
rect 15260 4162 15316 4172
rect 15484 4134 15540 4172
rect 15036 3948 15316 4004
rect 14924 2212 14980 2716
rect 15148 3668 15204 3678
rect 15148 3442 15204 3612
rect 15148 3390 15150 3442
rect 15202 3390 15204 3442
rect 15148 2772 15204 3390
rect 15260 2884 15316 3948
rect 15596 3556 15652 3566
rect 15596 3462 15652 3500
rect 15820 3220 15876 5740
rect 15820 3154 15876 3164
rect 15932 6468 15988 6478
rect 15932 5682 15988 6412
rect 16380 6468 16436 6860
rect 16604 6692 16660 6702
rect 16604 6598 16660 6636
rect 16156 6244 16212 6254
rect 16044 6132 16100 6142
rect 16044 6038 16100 6076
rect 15932 5630 15934 5682
rect 15986 5630 15988 5682
rect 15932 2996 15988 5630
rect 16156 5124 16212 6188
rect 16380 6020 16436 6412
rect 16380 5954 16436 5964
rect 16492 6466 16548 6478
rect 16492 6414 16494 6466
rect 16546 6414 16548 6466
rect 16380 5794 16436 5806
rect 16380 5742 16382 5794
rect 16434 5742 16436 5794
rect 16380 5682 16436 5742
rect 16380 5630 16382 5682
rect 16434 5630 16436 5682
rect 16380 5618 16436 5630
rect 16492 5348 16548 6414
rect 16716 5460 16772 7308
rect 16828 7298 16884 7308
rect 16828 6578 16884 6590
rect 16828 6526 16830 6578
rect 16882 6526 16884 6578
rect 16828 6020 16884 6526
rect 16828 5954 16884 5964
rect 17052 5908 17108 18620
rect 17500 18450 17556 18732
rect 17500 18398 17502 18450
rect 17554 18398 17556 18450
rect 17164 17554 17220 17566
rect 17164 17502 17166 17554
rect 17218 17502 17220 17554
rect 17164 14756 17220 17502
rect 17388 16996 17444 17006
rect 17164 14690 17220 14700
rect 17276 16324 17332 16334
rect 17276 15316 17332 16268
rect 17388 16212 17444 16940
rect 17388 16146 17444 16156
rect 17164 14084 17220 14094
rect 17164 10164 17220 14028
rect 17276 10276 17332 15260
rect 17388 14980 17444 14990
rect 17388 11954 17444 14924
rect 17388 11902 17390 11954
rect 17442 11902 17444 11954
rect 17388 11890 17444 11902
rect 17500 11508 17556 18398
rect 17612 17668 17668 19516
rect 17612 17602 17668 17612
rect 17724 19346 17780 19358
rect 17724 19294 17726 19346
rect 17778 19294 17780 19346
rect 17724 17108 17780 19294
rect 17836 19234 17892 19516
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 19170 17892 19182
rect 18060 19906 18116 19918
rect 18060 19854 18062 19906
rect 18114 19854 18116 19906
rect 18060 18674 18116 19854
rect 18060 18622 18062 18674
rect 18114 18622 18116 18674
rect 18060 18610 18116 18622
rect 18172 18900 18228 18910
rect 18172 18674 18228 18844
rect 18172 18622 18174 18674
rect 18226 18622 18228 18674
rect 18172 18610 18228 18622
rect 17836 18562 17892 18574
rect 17836 18510 17838 18562
rect 17890 18510 17892 18562
rect 17836 18340 17892 18510
rect 17948 18564 18004 18574
rect 17948 18470 18004 18508
rect 17836 18274 17892 18284
rect 18284 17780 18340 20748
rect 18396 20356 18452 22428
rect 18508 22146 18564 22158
rect 18508 22094 18510 22146
rect 18562 22094 18564 22146
rect 18508 21700 18564 22094
rect 18508 21634 18564 21644
rect 18508 21474 18564 21486
rect 18508 21422 18510 21474
rect 18562 21422 18564 21474
rect 18508 20468 18564 21422
rect 18620 21364 18676 23324
rect 18620 21298 18676 21308
rect 18732 21474 18788 21486
rect 18732 21422 18734 21474
rect 18786 21422 18788 21474
rect 18732 21028 18788 21422
rect 18732 20962 18788 20972
rect 18620 20580 18676 20590
rect 18620 20486 18676 20524
rect 18508 20402 18564 20412
rect 18396 20290 18452 20300
rect 18844 20244 18900 24892
rect 18620 20188 18900 20244
rect 18396 20132 18452 20142
rect 18396 20038 18452 20076
rect 18060 17724 18340 17780
rect 17948 17668 18004 17678
rect 17612 17052 17724 17108
rect 17612 15314 17668 17052
rect 17724 17014 17780 17052
rect 17836 17332 17892 17342
rect 17836 17106 17892 17276
rect 17836 17054 17838 17106
rect 17890 17054 17892 17106
rect 17836 17042 17892 17054
rect 17948 16660 18004 17612
rect 17612 15262 17614 15314
rect 17666 15262 17668 15314
rect 17612 15250 17668 15262
rect 17836 16604 18004 16660
rect 17836 13748 17892 16604
rect 17948 15876 18004 15886
rect 17948 15314 18004 15820
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 17948 15250 18004 15262
rect 18060 13748 18116 17724
rect 18284 17666 18340 17724
rect 18284 17614 18286 17666
rect 18338 17614 18340 17666
rect 18284 17602 18340 17614
rect 18620 17668 18676 20188
rect 18732 20018 18788 20030
rect 18732 19966 18734 20018
rect 18786 19966 18788 20018
rect 18732 18788 18788 19966
rect 18844 19460 18900 19470
rect 18844 19234 18900 19404
rect 18844 19182 18846 19234
rect 18898 19182 18900 19234
rect 18844 19170 18900 19182
rect 18732 18722 18788 18732
rect 18620 17574 18676 17612
rect 18844 18338 18900 18350
rect 18844 18286 18846 18338
rect 18898 18286 18900 18338
rect 18844 17668 18900 18286
rect 18172 17554 18228 17566
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 18172 17108 18228 17502
rect 18844 17220 18900 17612
rect 18844 17154 18900 17164
rect 18956 17332 19012 26852
rect 19180 24836 19236 27582
rect 21084 27300 21140 27310
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20076 26290 20132 26302
rect 20076 26238 20078 26290
rect 20130 26238 20132 26290
rect 19628 26178 19684 26190
rect 19628 26126 19630 26178
rect 19682 26126 19684 26178
rect 19628 25620 19684 26126
rect 19628 25554 19684 25564
rect 19404 25282 19460 25294
rect 19404 25230 19406 25282
rect 19458 25230 19460 25282
rect 19180 24770 19236 24780
rect 19292 24836 19348 24846
rect 19404 24836 19460 25230
rect 20076 25284 20132 26238
rect 20412 26178 20468 26190
rect 20412 26126 20414 26178
rect 20466 26126 20468 26178
rect 20300 25620 20356 25630
rect 20300 25526 20356 25564
rect 20412 25618 20468 26126
rect 20412 25566 20414 25618
rect 20466 25566 20468 25618
rect 20412 25554 20468 25566
rect 20636 25956 20692 25966
rect 20636 25506 20692 25900
rect 20636 25454 20638 25506
rect 20690 25454 20692 25506
rect 20636 25442 20692 25454
rect 20076 25228 20244 25284
rect 20188 25172 20244 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20188 25106 20244 25116
rect 19836 25050 20100 25060
rect 20860 24948 20916 24958
rect 20860 24854 20916 24892
rect 19292 24834 19460 24836
rect 19292 24782 19294 24834
rect 19346 24782 19460 24834
rect 19292 24780 19460 24782
rect 20972 24836 21028 24846
rect 19292 24770 19348 24780
rect 19852 24722 19908 24734
rect 19852 24670 19854 24722
rect 19906 24670 19908 24722
rect 19068 24612 19124 24622
rect 19516 24612 19572 24622
rect 19124 24556 19460 24612
rect 19068 24518 19124 24556
rect 19404 24164 19460 24556
rect 19516 24610 19684 24612
rect 19516 24558 19518 24610
rect 19570 24558 19684 24610
rect 19516 24556 19684 24558
rect 19516 24546 19572 24556
rect 19516 24164 19572 24174
rect 19404 24162 19572 24164
rect 19404 24110 19518 24162
rect 19570 24110 19572 24162
rect 19404 24108 19572 24110
rect 19516 24098 19572 24108
rect 19292 24052 19348 24062
rect 19292 23940 19348 23996
rect 19628 23940 19684 24556
rect 19292 23938 19684 23940
rect 19292 23886 19294 23938
rect 19346 23886 19684 23938
rect 19292 23884 19684 23886
rect 19852 23940 19908 24670
rect 20412 24612 20468 24622
rect 20412 24518 20468 24556
rect 19292 23874 19348 23884
rect 19852 23874 19908 23884
rect 19852 23716 19908 23726
rect 19852 23714 20244 23716
rect 19852 23662 19854 23714
rect 19906 23662 20244 23714
rect 19852 23660 20244 23662
rect 19852 23650 19908 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19852 23154 19908 23166
rect 19852 23102 19854 23154
rect 19906 23102 19908 23154
rect 19068 23042 19124 23054
rect 19068 22990 19070 23042
rect 19122 22990 19124 23042
rect 19068 22372 19124 22990
rect 19516 23042 19572 23054
rect 19516 22990 19518 23042
rect 19570 22990 19572 23042
rect 19068 22306 19124 22316
rect 19292 22370 19348 22382
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 22260 19348 22318
rect 19292 21810 19348 22204
rect 19292 21758 19294 21810
rect 19346 21758 19348 21810
rect 19292 21746 19348 21758
rect 19404 21700 19460 21710
rect 19180 20802 19236 20814
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 19180 20580 19236 20750
rect 19180 20244 19236 20524
rect 19180 20178 19236 20188
rect 19068 20130 19124 20142
rect 19068 20078 19070 20130
rect 19122 20078 19124 20130
rect 19068 19684 19124 20078
rect 19068 19618 19124 19628
rect 18172 17052 18676 17108
rect 18172 16882 18228 17052
rect 18172 16830 18174 16882
rect 18226 16830 18228 16882
rect 18172 16818 18228 16830
rect 18284 16884 18340 16894
rect 18172 16212 18228 16222
rect 18172 16098 18228 16156
rect 18172 16046 18174 16098
rect 18226 16046 18228 16098
rect 18172 16034 18228 16046
rect 18284 15876 18340 16828
rect 18284 15810 18340 15820
rect 18396 15986 18452 15998
rect 18396 15934 18398 15986
rect 18450 15934 18452 15986
rect 18396 14756 18452 15934
rect 18508 15652 18564 15662
rect 18508 15314 18564 15596
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 15250 18564 15262
rect 18620 15202 18676 17052
rect 18956 16882 19012 17276
rect 18956 16830 18958 16882
rect 19010 16830 19012 16882
rect 18956 16818 19012 16830
rect 19068 19460 19124 19470
rect 19068 18450 19124 19404
rect 19292 19122 19348 19134
rect 19292 19070 19294 19122
rect 19346 19070 19348 19122
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 16100 19124 18398
rect 19180 18562 19236 18574
rect 19180 18510 19182 18562
rect 19234 18510 19236 18562
rect 19180 16660 19236 18510
rect 19292 18004 19348 19070
rect 19292 17938 19348 17948
rect 19180 16594 19236 16604
rect 19180 16100 19236 16110
rect 19068 16098 19236 16100
rect 19068 16046 19182 16098
rect 19234 16046 19236 16098
rect 19068 16044 19236 16046
rect 19404 16100 19460 21644
rect 19516 20130 19572 22990
rect 19852 22148 19908 23102
rect 20188 23156 20244 23660
rect 20524 23714 20580 23726
rect 20524 23662 20526 23714
rect 20578 23662 20580 23714
rect 20300 23156 20356 23166
rect 20188 23100 20300 23156
rect 20524 23156 20580 23662
rect 20972 23716 21028 24780
rect 20972 23378 21028 23660
rect 20972 23326 20974 23378
rect 21026 23326 21028 23378
rect 20972 23314 21028 23326
rect 20636 23156 20692 23166
rect 20524 23154 20692 23156
rect 20524 23102 20638 23154
rect 20690 23102 20692 23154
rect 20524 23100 20692 23102
rect 20300 23062 20356 23100
rect 20076 22708 20132 22718
rect 20076 22482 20132 22652
rect 20076 22430 20078 22482
rect 20130 22430 20132 22482
rect 20076 22418 20132 22430
rect 19628 22092 19908 22148
rect 20524 22372 20580 22382
rect 20524 22258 20580 22316
rect 20524 22206 20526 22258
rect 20578 22206 20580 22258
rect 19628 21586 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21534 19630 21586
rect 19682 21534 19684 21586
rect 19628 21364 19684 21534
rect 19628 21298 19684 21308
rect 20524 21140 20580 22206
rect 20300 21084 20580 21140
rect 19740 20692 19796 20702
rect 19740 20580 19796 20636
rect 19628 20524 19796 20580
rect 19628 20468 19684 20524
rect 19628 20402 19684 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19516 20078 19518 20130
rect 19570 20078 19572 20130
rect 19516 20066 19572 20078
rect 19740 20018 19796 20030
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 19740 19458 19796 19966
rect 19740 19406 19742 19458
rect 19794 19406 19796 19458
rect 19740 19394 19796 19406
rect 20076 19346 20132 19358
rect 20076 19294 20078 19346
rect 20130 19294 20132 19346
rect 19740 19234 19796 19246
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19740 19124 19796 19182
rect 20076 19236 20132 19294
rect 20076 19170 20132 19180
rect 19740 19058 19796 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20300 18452 20356 21084
rect 20636 21028 20692 23100
rect 20860 22372 20916 22382
rect 20748 21700 20804 21710
rect 20748 21606 20804 21644
rect 20524 20972 20692 21028
rect 20524 20804 20580 20972
rect 20524 20738 20580 20748
rect 20636 20802 20692 20814
rect 20636 20750 20638 20802
rect 20690 20750 20692 20802
rect 20412 20690 20468 20702
rect 20412 20638 20414 20690
rect 20466 20638 20468 20690
rect 20412 19124 20468 20638
rect 20412 19058 20468 19068
rect 20636 19908 20692 20750
rect 20748 20690 20804 20702
rect 20748 20638 20750 20690
rect 20802 20638 20804 20690
rect 20748 20020 20804 20638
rect 20748 19954 20804 19964
rect 20412 18452 20468 18462
rect 20300 18396 20412 18452
rect 20188 18004 20244 18014
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19852 16882 19908 17052
rect 19852 16830 19854 16882
rect 19906 16830 19908 16882
rect 19852 16818 19908 16830
rect 20076 16324 20132 16334
rect 20076 16230 20132 16268
rect 19964 16100 20020 16110
rect 19404 16044 19684 16100
rect 19180 16034 19236 16044
rect 18620 15150 18622 15202
rect 18674 15150 18676 15202
rect 18620 15138 18676 15150
rect 18844 15988 18900 15998
rect 18844 15874 18900 15932
rect 18844 15822 18846 15874
rect 18898 15822 18900 15874
rect 18732 15092 18788 15102
rect 18732 14998 18788 15036
rect 18172 14644 18228 14654
rect 18172 13858 18228 14588
rect 18396 13972 18452 14700
rect 18396 13906 18452 13916
rect 18732 14756 18788 14766
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13794 18228 13806
rect 17836 13746 18004 13748
rect 17836 13694 17838 13746
rect 17890 13694 18004 13746
rect 17836 13692 18004 13694
rect 17836 13682 17892 13692
rect 17612 12962 17668 12974
rect 17612 12910 17614 12962
rect 17666 12910 17668 12962
rect 17612 12404 17668 12910
rect 17948 12404 18004 13692
rect 18060 13682 18116 13692
rect 18172 13636 18228 13646
rect 17948 12348 18116 12404
rect 17612 12338 17668 12348
rect 17724 12066 17780 12078
rect 17724 12014 17726 12066
rect 17778 12014 17780 12066
rect 17724 11954 17780 12014
rect 17724 11902 17726 11954
rect 17778 11902 17780 11954
rect 17724 11890 17780 11902
rect 18060 11788 18116 12348
rect 17836 11732 18116 11788
rect 17836 11666 17892 11676
rect 17500 11452 17892 11508
rect 17612 11282 17668 11294
rect 17612 11230 17614 11282
rect 17666 11230 17668 11282
rect 17612 10948 17668 11230
rect 17612 10882 17668 10892
rect 17724 10836 17780 10846
rect 17724 10742 17780 10780
rect 17276 10220 17668 10276
rect 17164 10108 17556 10164
rect 17388 9828 17444 9838
rect 17388 9734 17444 9772
rect 17164 9714 17220 9726
rect 17164 9662 17166 9714
rect 17218 9662 17220 9714
rect 17164 9492 17220 9662
rect 17164 9156 17220 9436
rect 17164 9090 17220 9100
rect 17500 8372 17556 10108
rect 17612 9266 17668 10220
rect 17612 9214 17614 9266
rect 17666 9214 17668 9266
rect 17612 9202 17668 9214
rect 17724 9714 17780 9726
rect 17724 9662 17726 9714
rect 17778 9662 17780 9714
rect 17276 7812 17332 7822
rect 17276 7476 17332 7756
rect 17500 7700 17556 8316
rect 17724 8258 17780 9662
rect 17836 9156 17892 11452
rect 18060 11172 18116 11182
rect 18060 11078 18116 11116
rect 18172 10836 18228 13580
rect 18732 13636 18788 14700
rect 18844 14530 18900 15822
rect 19628 15876 19684 16044
rect 19964 16006 20020 16044
rect 19628 15540 19684 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15484 19796 15540
rect 18844 14478 18846 14530
rect 18898 14478 18900 14530
rect 18844 14466 18900 14478
rect 18956 15428 19012 15438
rect 18732 13634 18900 13636
rect 18732 13582 18734 13634
rect 18786 13582 18900 13634
rect 18732 13580 18900 13582
rect 18732 13570 18788 13580
rect 18732 13412 18788 13422
rect 18284 13186 18340 13198
rect 18284 13134 18286 13186
rect 18338 13134 18340 13186
rect 18284 12404 18340 13134
rect 18284 12338 18340 12348
rect 18620 12066 18676 12078
rect 18620 12014 18622 12066
rect 18674 12014 18676 12066
rect 18620 11284 18676 12014
rect 18620 10948 18676 11228
rect 18620 10882 18676 10892
rect 18172 10780 18340 10836
rect 17948 10612 18004 10622
rect 17948 10518 18004 10556
rect 18172 10610 18228 10622
rect 18172 10558 18174 10610
rect 18226 10558 18228 10610
rect 18060 10500 18116 10510
rect 18060 10406 18116 10444
rect 18172 9940 18228 10558
rect 17836 9062 17892 9100
rect 17948 9884 18228 9940
rect 17948 8932 18004 9884
rect 18172 9716 18228 9726
rect 18172 9622 18228 9660
rect 17724 8206 17726 8258
rect 17778 8206 17780 8258
rect 17724 8194 17780 8206
rect 17836 8876 18004 8932
rect 18172 8930 18228 8942
rect 18172 8878 18174 8930
rect 18226 8878 18228 8930
rect 17612 8036 17668 8046
rect 17836 8036 17892 8876
rect 18060 8820 18116 8830
rect 18060 8726 18116 8764
rect 18172 8708 18228 8878
rect 18172 8642 18228 8652
rect 17612 8034 17780 8036
rect 17612 7982 17614 8034
rect 17666 7982 17780 8034
rect 17612 7980 17780 7982
rect 17612 7970 17668 7980
rect 17612 7700 17668 7710
rect 17500 7698 17668 7700
rect 17500 7646 17614 7698
rect 17666 7646 17668 7698
rect 17500 7644 17668 7646
rect 17276 7474 17444 7476
rect 17276 7422 17278 7474
rect 17330 7422 17444 7474
rect 17276 7420 17444 7422
rect 17276 7410 17332 7420
rect 16940 5852 17108 5908
rect 16828 5796 16884 5806
rect 16940 5796 16996 5852
rect 16828 5794 16996 5796
rect 16828 5742 16830 5794
rect 16882 5742 16996 5794
rect 16828 5740 16996 5742
rect 16828 5730 16884 5740
rect 16716 5404 16884 5460
rect 16492 5282 16548 5292
rect 16716 5236 16772 5246
rect 16716 5142 16772 5180
rect 16268 5124 16324 5134
rect 16156 5122 16324 5124
rect 16156 5070 16270 5122
rect 16322 5070 16324 5122
rect 16156 5068 16324 5070
rect 16268 5058 16324 5068
rect 16604 5122 16660 5134
rect 16604 5070 16606 5122
rect 16658 5070 16660 5122
rect 16044 4564 16100 4574
rect 16044 4470 16100 4508
rect 16604 4564 16660 5070
rect 16828 5012 16884 5404
rect 16940 5348 16996 5358
rect 16940 5254 16996 5292
rect 16604 4498 16660 4508
rect 16716 4956 16884 5012
rect 16268 4340 16324 4350
rect 16268 4246 16324 4284
rect 16716 4226 16772 4956
rect 16716 4174 16718 4226
rect 16770 4174 16772 4226
rect 16716 4162 16772 4174
rect 16492 3892 16548 3902
rect 16044 3668 16100 3678
rect 16044 3574 16100 3612
rect 16492 3666 16548 3836
rect 17052 3780 17108 5852
rect 17276 6020 17332 6030
rect 17052 3714 17108 3724
rect 17164 4340 17220 4350
rect 16492 3614 16494 3666
rect 16546 3614 16548 3666
rect 16492 3602 16548 3614
rect 17164 3554 17220 4284
rect 17164 3502 17166 3554
rect 17218 3502 17220 3554
rect 17164 3490 17220 3502
rect 17276 3108 17332 5964
rect 17388 5906 17444 7420
rect 17500 6916 17556 7644
rect 17612 7634 17668 7644
rect 17500 6850 17556 6860
rect 17388 5854 17390 5906
rect 17442 5854 17444 5906
rect 17388 5842 17444 5854
rect 17500 6690 17556 6702
rect 17500 6638 17502 6690
rect 17554 6638 17556 6690
rect 17500 5908 17556 6638
rect 17500 5842 17556 5852
rect 17612 5794 17668 5806
rect 17612 5742 17614 5794
rect 17666 5742 17668 5794
rect 17500 5010 17556 5022
rect 17500 4958 17502 5010
rect 17554 4958 17556 5010
rect 17500 3388 17556 4958
rect 17612 4450 17668 5742
rect 17724 5684 17780 7980
rect 17836 7970 17892 7980
rect 17948 8260 18004 8270
rect 17948 7698 18004 8204
rect 18284 8148 18340 10780
rect 18620 10610 18676 10622
rect 18620 10558 18622 10610
rect 18674 10558 18676 10610
rect 18620 10500 18676 10558
rect 18396 10444 18676 10500
rect 18396 9492 18452 10444
rect 18620 10276 18676 10286
rect 18396 9426 18452 9436
rect 18508 9826 18564 9838
rect 18508 9774 18510 9826
rect 18562 9774 18564 9826
rect 18508 8260 18564 9774
rect 18620 9716 18676 10220
rect 18620 9650 18676 9660
rect 18508 8194 18564 8204
rect 18732 8258 18788 13356
rect 18844 11396 18900 13580
rect 18956 11732 19012 15372
rect 19628 15314 19684 15326
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19404 15092 19460 15102
rect 19292 14644 19348 14654
rect 19068 12962 19124 12974
rect 19068 12910 19070 12962
rect 19122 12910 19124 12962
rect 19068 12740 19124 12910
rect 19068 12674 19124 12684
rect 19068 12516 19124 12526
rect 19068 12178 19124 12460
rect 19068 12126 19070 12178
rect 19122 12126 19124 12178
rect 19068 12114 19124 12126
rect 19180 12180 19236 12190
rect 18956 11666 19012 11676
rect 19068 11508 19124 11518
rect 19068 11414 19124 11452
rect 18844 11330 18900 11340
rect 19180 11394 19236 12124
rect 19292 11508 19348 14588
rect 19404 14530 19460 15036
rect 19404 14478 19406 14530
rect 19458 14478 19460 14530
rect 19404 14466 19460 14478
rect 19628 13972 19684 15262
rect 19740 14530 19796 15484
rect 19852 15426 19908 15438
rect 19852 15374 19854 15426
rect 19906 15374 19908 15426
rect 19852 15092 19908 15374
rect 19964 15316 20020 15326
rect 19964 15222 20020 15260
rect 19852 14756 19908 15036
rect 20188 14868 20244 17948
rect 20412 17668 20468 18396
rect 20300 17666 20468 17668
rect 20300 17614 20414 17666
rect 20466 17614 20468 17666
rect 20300 17612 20468 17614
rect 20300 17332 20356 17612
rect 20412 17602 20468 17612
rect 20524 18340 20580 18350
rect 20524 17444 20580 18284
rect 20636 17892 20692 19852
rect 20748 19012 20804 19022
rect 20748 18918 20804 18956
rect 20748 18452 20804 18462
rect 20748 18358 20804 18396
rect 20636 17826 20692 17836
rect 20300 17266 20356 17276
rect 20412 17388 20580 17444
rect 20748 17442 20804 17454
rect 20748 17390 20750 17442
rect 20802 17390 20804 17442
rect 20300 16884 20356 16894
rect 20300 16790 20356 16828
rect 20412 15426 20468 17388
rect 20748 17220 20804 17390
rect 20748 17154 20804 17164
rect 20524 16436 20580 16446
rect 20524 16098 20580 16380
rect 20860 16436 20916 22316
rect 21084 20242 21140 27244
rect 21644 26628 21700 26638
rect 21196 26404 21252 26414
rect 21196 26310 21252 26348
rect 21644 26290 21700 26572
rect 21644 26238 21646 26290
rect 21698 26238 21700 26290
rect 21644 26226 21700 26238
rect 21756 26292 21812 27692
rect 22764 27076 22820 27086
rect 22764 26982 22820 27020
rect 22652 26962 22708 26974
rect 22652 26910 22654 26962
rect 22706 26910 22708 26962
rect 22652 26908 22708 26910
rect 22540 26852 22708 26908
rect 22876 26852 22932 26862
rect 22540 26402 22596 26852
rect 22876 26758 22932 26796
rect 23100 26516 23156 27916
rect 25228 27858 25284 27870
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 24220 27748 24276 27758
rect 24220 27654 24276 27692
rect 25228 27748 25284 27806
rect 25228 27682 25284 27692
rect 25676 27186 25732 28364
rect 25900 27636 25956 28700
rect 26572 28644 26628 30942
rect 26796 30994 27076 30996
rect 26796 30942 27022 30994
rect 27074 30942 27076 30994
rect 26796 30940 27076 30942
rect 26796 30434 26852 30940
rect 27020 30930 27076 30940
rect 26796 30382 26798 30434
rect 26850 30382 26852 30434
rect 26796 30370 26852 30382
rect 28588 30212 28644 31892
rect 29260 31890 29428 31892
rect 29260 31838 29374 31890
rect 29426 31838 29428 31890
rect 29260 31836 29428 31838
rect 29372 31826 29428 31836
rect 29596 31668 29652 31892
rect 29596 31602 29652 31612
rect 30156 31220 30212 31230
rect 30268 31220 30324 31892
rect 30156 31218 30324 31220
rect 30156 31166 30158 31218
rect 30210 31166 30324 31218
rect 30156 31164 30324 31166
rect 30156 31154 30212 31164
rect 28476 30156 28644 30212
rect 29372 31106 29428 31118
rect 29372 31054 29374 31106
rect 29426 31054 29428 31106
rect 26684 29988 26740 29998
rect 26684 29894 26740 29932
rect 28364 29426 28420 29438
rect 28364 29374 28366 29426
rect 28418 29374 28420 29426
rect 27916 29316 27972 29326
rect 27916 29222 27972 29260
rect 28364 29316 28420 29374
rect 28364 29250 28420 29260
rect 28476 28866 28532 30156
rect 28476 28814 28478 28866
rect 28530 28814 28532 28866
rect 28476 28802 28532 28814
rect 28588 29652 28644 29662
rect 27916 28644 27972 28654
rect 28588 28644 28644 29596
rect 26572 28578 26628 28588
rect 27804 28588 27916 28644
rect 27692 28532 27748 28542
rect 27692 28438 27748 28476
rect 26124 28420 26180 28430
rect 26012 28084 26068 28094
rect 26012 27990 26068 28028
rect 26124 27970 26180 28364
rect 26124 27918 26126 27970
rect 26178 27918 26180 27970
rect 26124 27906 26180 27918
rect 26684 28084 26740 28094
rect 26012 27636 26068 27646
rect 25900 27634 26068 27636
rect 25900 27582 26014 27634
rect 26066 27582 26068 27634
rect 25900 27580 26068 27582
rect 25676 27134 25678 27186
rect 25730 27134 25732 27186
rect 25676 27122 25732 27134
rect 22540 26350 22542 26402
rect 22594 26350 22596 26402
rect 22540 26338 22596 26350
rect 22764 26460 23156 26516
rect 23324 26962 23380 26974
rect 23324 26910 23326 26962
rect 23378 26910 23380 26962
rect 21756 26226 21812 26236
rect 22092 26178 22148 26190
rect 22092 26126 22094 26178
rect 22146 26126 22148 26178
rect 22092 26068 22148 26126
rect 22092 26002 22148 26012
rect 21420 25956 21476 25966
rect 21420 25618 21476 25900
rect 22540 25732 22596 25742
rect 22540 25638 22596 25676
rect 21420 25566 21422 25618
rect 21474 25566 21476 25618
rect 21420 25554 21476 25566
rect 22764 25620 22820 26460
rect 23324 26404 23380 26910
rect 23436 26962 23492 26974
rect 23436 26910 23438 26962
rect 23490 26910 23492 26962
rect 23436 26628 23492 26910
rect 23436 26562 23492 26572
rect 23548 26852 23604 26862
rect 23324 26348 23492 26404
rect 22988 26290 23044 26302
rect 22988 26238 22990 26290
rect 23042 26238 23044 26290
rect 22876 26180 22932 26190
rect 22876 25730 22932 26124
rect 22988 25844 23044 26238
rect 23324 26180 23380 26190
rect 22988 25778 23044 25788
rect 23100 26178 23380 26180
rect 23100 26126 23326 26178
rect 23378 26126 23380 26178
rect 23100 26124 23380 26126
rect 22876 25678 22878 25730
rect 22930 25678 22932 25730
rect 22876 25666 22932 25678
rect 22764 25508 22820 25564
rect 23100 25620 23156 26124
rect 23324 26114 23380 26124
rect 23436 26068 23492 26348
rect 23436 26002 23492 26012
rect 23100 25526 23156 25564
rect 22764 25452 23044 25508
rect 22988 24724 23044 25452
rect 23324 25060 23380 25070
rect 23100 24724 23156 24734
rect 22988 24722 23156 24724
rect 22988 24670 23102 24722
rect 23154 24670 23156 24722
rect 22988 24668 23156 24670
rect 23100 24658 23156 24668
rect 22876 24610 22932 24622
rect 22876 24558 22878 24610
rect 22930 24558 22932 24610
rect 22876 24500 22932 24558
rect 22876 24164 22932 24444
rect 23324 24500 23380 25004
rect 23548 24836 23604 26796
rect 23660 26852 23716 26862
rect 24332 26852 24388 26862
rect 23660 26850 23828 26852
rect 23660 26798 23662 26850
rect 23714 26798 23828 26850
rect 23660 26796 23828 26798
rect 23660 26786 23716 26796
rect 23772 26290 23828 26796
rect 23772 26238 23774 26290
rect 23826 26238 23828 26290
rect 23772 26226 23828 26238
rect 24220 26292 24276 26302
rect 24220 26198 24276 26236
rect 24332 26290 24388 26796
rect 24332 26238 24334 26290
rect 24386 26238 24388 26290
rect 24332 26226 24388 26238
rect 24780 26628 24836 26638
rect 23996 26180 24052 26190
rect 23996 26086 24052 26124
rect 23772 25844 23828 25854
rect 23772 25618 23828 25788
rect 23772 25566 23774 25618
rect 23826 25566 23828 25618
rect 23772 25554 23828 25566
rect 23884 25732 23940 25742
rect 23884 25172 23940 25676
rect 24668 25620 24724 25630
rect 24668 25526 24724 25564
rect 24780 25508 24836 26572
rect 25900 26290 25956 26302
rect 25900 26238 25902 26290
rect 25954 26238 25956 26290
rect 25900 26180 25956 26238
rect 25900 26114 25956 26124
rect 26012 26178 26068 27580
rect 26684 27186 26740 28028
rect 27132 28084 27188 28094
rect 27132 27858 27188 28028
rect 27692 28084 27748 28094
rect 27804 28084 27860 28588
rect 27916 28578 27972 28588
rect 28476 28588 28644 28644
rect 29148 28644 29204 28654
rect 27692 28082 27860 28084
rect 27692 28030 27694 28082
rect 27746 28030 27860 28082
rect 27692 28028 27860 28030
rect 28140 28532 28196 28542
rect 27692 28018 27748 28028
rect 27132 27806 27134 27858
rect 27186 27806 27188 27858
rect 27132 27794 27188 27806
rect 26908 27746 26964 27758
rect 26908 27694 26910 27746
rect 26962 27694 26964 27746
rect 26908 27524 26964 27694
rect 28140 27746 28196 28476
rect 28476 27858 28532 28588
rect 29148 28550 29204 28588
rect 29372 28532 29428 31054
rect 30156 30996 30212 31006
rect 29820 30210 29876 30222
rect 29820 30158 29822 30210
rect 29874 30158 29876 30210
rect 29820 29650 29876 30158
rect 29820 29598 29822 29650
rect 29874 29598 29876 29650
rect 29820 29586 29876 29598
rect 30044 29428 30100 29438
rect 29596 29426 30100 29428
rect 29596 29374 30046 29426
rect 30098 29374 30100 29426
rect 29596 29372 30100 29374
rect 29372 28466 29428 28476
rect 29484 28644 29540 28654
rect 29484 28530 29540 28588
rect 29484 28478 29486 28530
rect 29538 28478 29540 28530
rect 29484 28466 29540 28478
rect 29596 27970 29652 29372
rect 30044 29362 30100 29372
rect 29596 27918 29598 27970
rect 29650 27918 29652 27970
rect 29596 27906 29652 27918
rect 30044 28644 30100 28654
rect 30156 28644 30212 30940
rect 31500 30996 31556 33292
rect 31948 33236 32004 34972
rect 32396 35028 32452 35038
rect 34076 35028 34132 38220
rect 34300 38164 34356 38558
rect 34300 38098 34356 38108
rect 34524 38052 34580 38062
rect 34524 37958 34580 37996
rect 34636 37940 34692 37950
rect 34636 37846 34692 37884
rect 34300 37604 34356 37614
rect 34300 37490 34356 37548
rect 34300 37438 34302 37490
rect 34354 37438 34356 37490
rect 34300 37426 34356 37438
rect 34188 37266 34244 37278
rect 34412 37268 34468 37278
rect 34188 37214 34190 37266
rect 34242 37214 34244 37266
rect 34188 37156 34244 37214
rect 34188 37090 34244 37100
rect 34300 37212 34412 37268
rect 34300 36594 34356 37212
rect 34412 37174 34468 37212
rect 34748 37156 34804 38612
rect 34748 37062 34804 37100
rect 34860 38612 35028 38668
rect 36652 38668 36708 40684
rect 36876 39844 36932 39854
rect 36652 38612 36820 38668
rect 34860 36932 34916 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 38052 35140 38062
rect 35084 37958 35140 37996
rect 35196 38050 35252 38062
rect 35196 37998 35198 38050
rect 35250 37998 35252 38050
rect 34972 37938 35028 37950
rect 34972 37886 34974 37938
rect 35026 37886 35028 37938
rect 34972 37268 35028 37886
rect 35196 37492 35252 37998
rect 35420 38050 35476 38062
rect 35420 37998 35422 38050
rect 35474 37998 35476 38050
rect 35196 37436 35364 37492
rect 35196 37268 35252 37278
rect 34972 37212 35196 37268
rect 35196 37174 35252 37212
rect 34972 37044 35028 37054
rect 35308 37044 35364 37436
rect 35420 37156 35476 37998
rect 35644 37828 35700 37838
rect 35644 37490 35700 37772
rect 35644 37438 35646 37490
rect 35698 37438 35700 37490
rect 35644 37426 35700 37438
rect 35420 37090 35476 37100
rect 35756 37156 35812 37166
rect 35028 36988 35364 37044
rect 34972 36950 35028 36988
rect 34300 36542 34302 36594
rect 34354 36542 34356 36594
rect 34300 36530 34356 36542
rect 34748 36876 34916 36932
rect 35196 36876 35460 36886
rect 34636 36484 34692 36494
rect 34524 36370 34580 36382
rect 34524 36318 34526 36370
rect 34578 36318 34580 36370
rect 34188 36036 34244 36046
rect 34188 35922 34244 35980
rect 34188 35870 34190 35922
rect 34242 35870 34244 35922
rect 34188 35858 34244 35870
rect 34524 35924 34580 36318
rect 34524 35810 34580 35868
rect 34524 35758 34526 35810
rect 34578 35758 34580 35810
rect 34524 35746 34580 35758
rect 34636 35810 34692 36428
rect 34636 35758 34638 35810
rect 34690 35758 34692 35810
rect 34636 35476 34692 35758
rect 34636 35410 34692 35420
rect 34636 35028 34692 35038
rect 34076 35026 34692 35028
rect 34076 34974 34638 35026
rect 34690 34974 34692 35026
rect 34076 34972 34692 34974
rect 32396 34934 32452 34972
rect 32508 34804 32564 34814
rect 32508 34710 32564 34748
rect 34636 34692 34692 34972
rect 34636 34626 34692 34636
rect 33404 34356 33460 34366
rect 33404 34262 33460 34300
rect 33852 34356 33908 34366
rect 33852 34262 33908 34300
rect 33068 34242 33124 34254
rect 33068 34190 33070 34242
rect 33122 34190 33124 34242
rect 32172 34132 32228 34142
rect 32172 34038 32228 34076
rect 32172 33348 32228 33358
rect 32172 33254 32228 33292
rect 33068 33348 33124 34190
rect 34412 34132 34468 34142
rect 34748 34132 34804 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35644 36484 35700 36494
rect 35644 36390 35700 36428
rect 35532 36372 35588 36382
rect 34860 35924 34916 35934
rect 34860 35830 34916 35868
rect 35532 35922 35588 36316
rect 35532 35870 35534 35922
rect 35586 35870 35588 35922
rect 35532 35858 35588 35870
rect 35644 35924 35700 35934
rect 35644 35830 35700 35868
rect 34972 35812 35028 35822
rect 34972 35698 35028 35756
rect 34972 35646 34974 35698
rect 35026 35646 35028 35698
rect 34972 35634 35028 35646
rect 35420 35698 35476 35710
rect 35420 35646 35422 35698
rect 35474 35646 35476 35698
rect 35420 35476 35476 35646
rect 35756 35588 35812 37100
rect 36204 35924 36260 35934
rect 36204 35698 36260 35868
rect 36204 35646 36206 35698
rect 36258 35646 36260 35698
rect 36204 35634 36260 35646
rect 36428 35812 36484 35822
rect 36428 35698 36484 35756
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 36428 35634 36484 35646
rect 34972 35420 35476 35476
rect 35644 35532 35812 35588
rect 35980 35586 36036 35598
rect 35980 35534 35982 35586
rect 36034 35534 36036 35586
rect 34972 35140 35028 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34860 34692 34916 34702
rect 34972 34692 35028 35084
rect 34916 34636 35028 34692
rect 35084 34916 35140 34926
rect 34860 34598 34916 34636
rect 34972 34132 35028 34142
rect 34748 34130 35028 34132
rect 34748 34078 34974 34130
rect 35026 34078 35028 34130
rect 34748 34076 35028 34078
rect 34412 34038 34468 34076
rect 34972 34066 35028 34076
rect 35084 33572 35140 34860
rect 35532 34804 35588 34814
rect 35644 34804 35700 35532
rect 35980 35140 36036 35534
rect 36764 35252 36820 38612
rect 36876 37378 36932 39788
rect 36988 38164 37044 44044
rect 37324 42980 37380 44268
rect 37324 42914 37380 42924
rect 37548 43428 37604 43438
rect 37548 42866 37604 43372
rect 37660 43204 37716 47516
rect 37996 45444 38052 48302
rect 38556 48356 38612 48366
rect 38612 48300 38836 48356
rect 38556 48262 38612 48300
rect 38332 48244 38388 48254
rect 38780 48244 38836 48300
rect 38892 48244 38948 48254
rect 38780 48242 38948 48244
rect 38780 48190 38894 48242
rect 38946 48190 38948 48242
rect 38780 48188 38948 48190
rect 38332 48150 38388 48188
rect 38108 47348 38164 47358
rect 38108 47254 38164 47292
rect 38556 45780 38612 45790
rect 38556 45778 38724 45780
rect 38556 45726 38558 45778
rect 38610 45726 38724 45778
rect 38556 45724 38724 45726
rect 38556 45714 38612 45724
rect 38668 45556 38724 45724
rect 38892 45778 38948 48188
rect 38892 45726 38894 45778
rect 38946 45726 38948 45778
rect 38892 45714 38948 45726
rect 39004 45556 39060 48412
rect 39116 48244 39172 48254
rect 39340 48244 39396 50372
rect 39788 49924 39844 50652
rect 39900 50484 39956 50494
rect 39900 50390 39956 50428
rect 39900 49924 39956 49934
rect 39788 49922 39956 49924
rect 39788 49870 39902 49922
rect 39954 49870 39956 49922
rect 39788 49868 39956 49870
rect 39564 49812 39620 49822
rect 39452 49810 39620 49812
rect 39452 49758 39566 49810
rect 39618 49758 39620 49810
rect 39452 49756 39620 49758
rect 39452 49028 39508 49756
rect 39564 49746 39620 49756
rect 39564 49140 39620 49150
rect 39564 49046 39620 49084
rect 39452 48934 39508 48972
rect 39676 48466 39732 48478
rect 39676 48414 39678 48466
rect 39730 48414 39732 48466
rect 39452 48244 39508 48254
rect 39340 48188 39452 48244
rect 39116 47124 39172 48188
rect 39340 48018 39396 48030
rect 39340 47966 39342 48018
rect 39394 47966 39396 48018
rect 39340 47346 39396 47966
rect 39452 47460 39508 48188
rect 39676 47684 39732 48414
rect 39788 48356 39844 49868
rect 39900 49858 39956 49868
rect 40012 48580 40068 51324
rect 40908 51156 40964 51166
rect 41020 51156 41076 51324
rect 41132 51314 41188 51324
rect 41244 51938 41300 51950
rect 41244 51886 41246 51938
rect 41298 51886 41300 51938
rect 41244 51156 41300 51886
rect 42028 51492 42084 52110
rect 42252 52164 42308 52174
rect 42028 51378 42084 51436
rect 42028 51326 42030 51378
rect 42082 51326 42084 51378
rect 42028 51314 42084 51326
rect 42140 51716 42196 51726
rect 41020 51100 41300 51156
rect 40908 51062 40964 51100
rect 39788 48290 39844 48300
rect 39900 48524 40068 48580
rect 40236 49138 40292 49150
rect 40236 49086 40238 49138
rect 40290 49086 40292 49138
rect 40236 48580 40292 49086
rect 39788 47684 39844 47694
rect 39676 47682 39844 47684
rect 39676 47630 39790 47682
rect 39842 47630 39844 47682
rect 39676 47628 39844 47630
rect 39788 47618 39844 47628
rect 39564 47460 39620 47470
rect 39452 47458 39620 47460
rect 39452 47406 39566 47458
rect 39618 47406 39620 47458
rect 39452 47404 39620 47406
rect 39564 47394 39620 47404
rect 39900 47458 39956 48524
rect 40236 48514 40292 48524
rect 40012 48354 40068 48366
rect 40012 48302 40014 48354
rect 40066 48302 40068 48354
rect 40012 48244 40068 48302
rect 40012 48178 40068 48188
rect 40236 48242 40292 48254
rect 40236 48190 40238 48242
rect 40290 48190 40292 48242
rect 40236 48132 40292 48190
rect 39900 47406 39902 47458
rect 39954 47406 39956 47458
rect 39340 47294 39342 47346
rect 39394 47294 39396 47346
rect 39340 47236 39396 47294
rect 39340 47170 39396 47180
rect 39116 47058 39172 47068
rect 39900 46900 39956 47406
rect 40124 48020 40180 48030
rect 40124 47234 40180 47964
rect 40236 47572 40292 48076
rect 41020 48132 41076 48142
rect 41020 48038 41076 48076
rect 40236 47506 40292 47516
rect 40124 47182 40126 47234
rect 40178 47182 40180 47234
rect 40124 47170 40180 47182
rect 39900 46834 39956 46844
rect 40012 47124 40068 47134
rect 38668 45500 39060 45556
rect 39116 45890 39172 45902
rect 39116 45838 39118 45890
rect 39170 45838 39172 45890
rect 37996 45388 38164 45444
rect 37996 45220 38052 45230
rect 37996 45126 38052 45164
rect 37884 45108 37940 45118
rect 37884 45014 37940 45052
rect 38108 43764 38164 45388
rect 38220 45108 38276 45118
rect 38556 45108 38612 45118
rect 38220 45106 38612 45108
rect 38220 45054 38222 45106
rect 38274 45054 38558 45106
rect 38610 45054 38612 45106
rect 38220 45052 38612 45054
rect 38220 45042 38276 45052
rect 38556 45042 38612 45052
rect 38668 44436 38724 45500
rect 38780 45106 38836 45118
rect 38780 45054 38782 45106
rect 38834 45054 38836 45106
rect 38780 44772 38836 45054
rect 38780 44706 38836 44716
rect 39116 44884 39172 45838
rect 39452 45780 39508 45790
rect 39452 45686 39508 45724
rect 40012 45330 40068 47068
rect 41020 46900 41076 46910
rect 41020 46806 41076 46844
rect 40012 45278 40014 45330
rect 40066 45278 40068 45330
rect 40012 45266 40068 45278
rect 40124 45666 40180 45678
rect 40124 45614 40126 45666
rect 40178 45614 40180 45666
rect 39452 45108 39508 45118
rect 39452 45014 39508 45052
rect 39788 45106 39844 45118
rect 39788 45054 39790 45106
rect 39842 45054 39844 45106
rect 38668 44322 38724 44380
rect 39116 44434 39172 44828
rect 39788 44996 39844 45054
rect 39116 44382 39118 44434
rect 39170 44382 39172 44434
rect 39116 44370 39172 44382
rect 39676 44436 39732 44446
rect 39676 44342 39732 44380
rect 38668 44270 38670 44322
rect 38722 44270 38724 44322
rect 38332 44098 38388 44110
rect 38332 44046 38334 44098
rect 38386 44046 38388 44098
rect 38332 43876 38388 44046
rect 38332 43810 38388 43820
rect 38108 43708 38276 43764
rect 38108 43540 38164 43550
rect 38108 43446 38164 43484
rect 37884 43428 37940 43438
rect 37884 43334 37940 43372
rect 37660 43148 38052 43204
rect 37548 42814 37550 42866
rect 37602 42814 37604 42866
rect 37548 42802 37604 42814
rect 37884 42980 37940 42990
rect 37772 40404 37828 40414
rect 37548 40402 37828 40404
rect 37548 40350 37774 40402
rect 37826 40350 37828 40402
rect 37548 40348 37828 40350
rect 37548 39842 37604 40348
rect 37772 40338 37828 40348
rect 37548 39790 37550 39842
rect 37602 39790 37604 39842
rect 37212 39618 37268 39630
rect 37212 39566 37214 39618
rect 37266 39566 37268 39618
rect 37212 39508 37268 39566
rect 37212 39442 37268 39452
rect 37436 39508 37492 39518
rect 37436 39414 37492 39452
rect 37548 38274 37604 39790
rect 37548 38222 37550 38274
rect 37602 38222 37604 38274
rect 37548 38210 37604 38222
rect 37772 38276 37828 38286
rect 37884 38276 37940 42924
rect 37996 39508 38052 43148
rect 38108 42868 38164 42878
rect 38220 42868 38276 43708
rect 38668 43428 38724 44270
rect 38780 44324 38836 44334
rect 38780 43650 38836 44268
rect 39228 44212 39284 44222
rect 39228 44118 39284 44156
rect 38780 43598 38782 43650
rect 38834 43598 38836 43650
rect 38780 43586 38836 43598
rect 39004 44098 39060 44110
rect 39004 44046 39006 44098
rect 39058 44046 39060 44098
rect 39004 43652 39060 44046
rect 39788 43652 39844 44940
rect 40124 44882 40180 45614
rect 40124 44830 40126 44882
rect 40178 44830 40180 44882
rect 40124 44212 40180 44830
rect 40460 45666 40516 45678
rect 40460 45614 40462 45666
rect 40514 45614 40516 45666
rect 40460 44436 40516 45614
rect 41244 45332 41300 51100
rect 42140 50818 42196 51660
rect 42252 51266 42308 52108
rect 42588 52164 42644 54236
rect 42924 53730 42980 55132
rect 44828 55188 44884 55198
rect 45388 55188 45444 55198
rect 44828 55094 44884 55132
rect 45276 55186 45444 55188
rect 45276 55134 45390 55186
rect 45442 55134 45444 55186
rect 45276 55132 45444 55134
rect 44940 55076 44996 55086
rect 44940 54852 44996 55020
rect 45164 55076 45220 55086
rect 45164 54982 45220 55020
rect 44716 54796 44996 54852
rect 44716 54626 44772 54796
rect 45052 54740 45108 54750
rect 45276 54740 45332 55132
rect 45388 55122 45444 55132
rect 45500 55188 45556 55198
rect 45500 55094 45556 55132
rect 45724 55188 45780 55198
rect 45724 55094 45780 55132
rect 46844 55186 46900 55198
rect 46844 55134 46846 55186
rect 46898 55134 46900 55186
rect 45052 54738 45332 54740
rect 45052 54686 45054 54738
rect 45106 54686 45332 54738
rect 45052 54684 45332 54686
rect 45052 54674 45108 54684
rect 44716 54574 44718 54626
rect 44770 54574 44772 54626
rect 44716 54562 44772 54574
rect 44828 54626 44884 54638
rect 44828 54574 44830 54626
rect 44882 54574 44884 54626
rect 43484 54516 43540 54526
rect 44380 54516 44436 54526
rect 43540 54460 43764 54516
rect 43484 54422 43540 54460
rect 42924 53678 42926 53730
rect 42978 53678 42980 53730
rect 42924 53666 42980 53678
rect 43596 53844 43652 53854
rect 43596 53618 43652 53788
rect 43596 53566 43598 53618
rect 43650 53566 43652 53618
rect 43596 52386 43652 53566
rect 43708 53618 43764 54460
rect 44380 54422 44436 54460
rect 43820 54402 43876 54414
rect 43820 54350 43822 54402
rect 43874 54350 43876 54402
rect 43820 53844 43876 54350
rect 43820 53778 43876 53788
rect 43708 53566 43710 53618
rect 43762 53566 43764 53618
rect 43708 53554 43764 53566
rect 43932 53620 43988 53630
rect 43932 53526 43988 53564
rect 44828 53620 44884 54574
rect 46844 54628 46900 55134
rect 46844 54534 46900 54572
rect 46956 55186 47012 55198
rect 46956 55134 46958 55186
rect 47010 55134 47012 55186
rect 46396 54514 46452 54526
rect 46396 54462 46398 54514
rect 46450 54462 46452 54514
rect 46172 54402 46228 54414
rect 46172 54350 46174 54402
rect 46226 54350 46228 54402
rect 46172 53956 46228 54350
rect 46172 53862 46228 53900
rect 44828 53554 44884 53564
rect 43596 52334 43598 52386
rect 43650 52334 43652 52386
rect 43596 52322 43652 52334
rect 46396 53506 46452 54462
rect 46956 54180 47012 55134
rect 47068 55188 47124 55198
rect 47068 54514 47124 55132
rect 47516 55188 47572 55198
rect 47852 55188 47908 55198
rect 47516 55186 47908 55188
rect 47516 55134 47518 55186
rect 47570 55134 47854 55186
rect 47906 55134 47908 55186
rect 47516 55132 47908 55134
rect 47516 55122 47572 55132
rect 47852 55122 47908 55132
rect 48076 55076 48132 55086
rect 47964 55074 48132 55076
rect 47964 55022 48078 55074
rect 48130 55022 48132 55074
rect 47964 55020 48132 55022
rect 47964 54852 48020 55020
rect 48076 55010 48132 55020
rect 47068 54462 47070 54514
rect 47122 54462 47124 54514
rect 47068 54450 47124 54462
rect 47404 54796 48020 54852
rect 47404 54738 47460 54796
rect 47404 54686 47406 54738
rect 47458 54686 47460 54738
rect 46956 54114 47012 54124
rect 47292 53956 47348 53966
rect 47404 53956 47460 54686
rect 47628 54628 47684 54638
rect 47516 54514 47572 54526
rect 47516 54462 47518 54514
rect 47570 54462 47572 54514
rect 47516 54180 47572 54462
rect 47628 54514 47684 54572
rect 47628 54462 47630 54514
rect 47682 54462 47684 54514
rect 47628 54450 47684 54462
rect 47516 54114 47572 54124
rect 47292 53954 47460 53956
rect 47292 53902 47294 53954
rect 47346 53902 47460 53954
rect 47292 53900 47460 53902
rect 47292 53890 47348 53900
rect 46508 53844 46564 53854
rect 46508 53842 47012 53844
rect 46508 53790 46510 53842
rect 46562 53790 47012 53842
rect 46508 53788 47012 53790
rect 46508 53778 46564 53788
rect 46956 53732 47012 53788
rect 47180 53732 47236 53742
rect 46956 53730 47124 53732
rect 46956 53678 46958 53730
rect 47010 53678 47124 53730
rect 46956 53676 47124 53678
rect 46956 53666 47012 53676
rect 46396 53454 46398 53506
rect 46450 53454 46452 53506
rect 43260 52274 43316 52286
rect 43260 52222 43262 52274
rect 43314 52222 43316 52274
rect 42588 52098 42644 52108
rect 43148 52162 43204 52174
rect 43148 52110 43150 52162
rect 43202 52110 43204 52162
rect 43148 51716 43204 52110
rect 43148 51650 43204 51660
rect 42700 51492 42756 51502
rect 43260 51492 43316 52222
rect 42700 51490 43316 51492
rect 42700 51438 42702 51490
rect 42754 51438 43316 51490
rect 42700 51436 43316 51438
rect 42700 51426 42756 51436
rect 42252 51214 42254 51266
rect 42306 51214 42308 51266
rect 42252 51202 42308 51214
rect 43260 51266 43316 51436
rect 43484 52162 43540 52174
rect 43484 52110 43486 52162
rect 43538 52110 43540 52162
rect 43260 51214 43262 51266
rect 43314 51214 43316 51266
rect 43260 51202 43316 51214
rect 43372 51378 43428 51390
rect 43372 51326 43374 51378
rect 43426 51326 43428 51378
rect 43372 50932 43428 51326
rect 42140 50766 42142 50818
rect 42194 50766 42196 50818
rect 42140 50754 42196 50766
rect 42476 50876 43428 50932
rect 42476 50818 42532 50876
rect 42476 50766 42478 50818
rect 42530 50766 42532 50818
rect 42476 50754 42532 50766
rect 42476 50596 42532 50606
rect 42476 50502 42532 50540
rect 43484 50596 43540 52110
rect 43932 52164 43988 52174
rect 43932 50596 43988 52108
rect 44940 52164 44996 52174
rect 44044 51268 44100 51278
rect 44044 51174 44100 51212
rect 44268 50932 44324 50942
rect 44044 50596 44100 50606
rect 43932 50594 44100 50596
rect 43932 50542 44046 50594
rect 44098 50542 44100 50594
rect 43932 50540 44100 50542
rect 43484 50530 43540 50540
rect 44044 50530 44100 50540
rect 44156 50484 44212 50494
rect 44156 50390 44212 50428
rect 43036 49924 43092 49934
rect 43036 49830 43092 49868
rect 43148 49922 43204 49934
rect 43148 49870 43150 49922
rect 43202 49870 43204 49922
rect 43148 49364 43204 49870
rect 43372 49812 43428 49822
rect 43372 49718 43428 49756
rect 43148 49308 43428 49364
rect 42252 49028 42308 49038
rect 42812 49028 42868 49038
rect 42252 48934 42308 48972
rect 42364 48972 42812 49028
rect 42364 48466 42420 48972
rect 42812 48934 42868 48972
rect 43260 49028 43316 49038
rect 43260 48934 43316 48972
rect 42924 48916 42980 48926
rect 42924 48822 42980 48860
rect 42364 48414 42366 48466
rect 42418 48414 42420 48466
rect 42364 48402 42420 48414
rect 43036 48804 43092 48814
rect 42140 48356 42196 48366
rect 42140 48262 42196 48300
rect 42476 48356 42532 48366
rect 42476 48262 42532 48300
rect 42588 48242 42644 48254
rect 42588 48190 42590 48242
rect 42642 48190 42644 48242
rect 42588 47348 42644 48190
rect 42140 47292 42644 47348
rect 42028 46788 42084 46798
rect 41244 45266 41300 45276
rect 41356 46674 41412 46686
rect 41356 46622 41358 46674
rect 41410 46622 41412 46674
rect 40460 44370 40516 44380
rect 40908 45220 40964 45230
rect 40908 44996 40964 45164
rect 41244 45106 41300 45118
rect 41244 45054 41246 45106
rect 41298 45054 41300 45106
rect 41020 44996 41076 45006
rect 40908 44994 41076 44996
rect 40908 44942 41022 44994
rect 41074 44942 41076 44994
rect 40908 44940 41076 44942
rect 40124 44146 40180 44156
rect 39004 43596 39844 43652
rect 38668 43372 38836 43428
rect 38668 42980 38724 42990
rect 38108 42866 38500 42868
rect 38108 42814 38110 42866
rect 38162 42814 38500 42866
rect 38108 42812 38500 42814
rect 38108 42802 38164 42812
rect 38220 39732 38276 42812
rect 38444 42754 38500 42812
rect 38444 42702 38446 42754
rect 38498 42702 38500 42754
rect 38444 42690 38500 42702
rect 38556 42756 38612 42766
rect 38556 42662 38612 42700
rect 38668 42196 38724 42924
rect 38668 42102 38724 42140
rect 38780 41748 38836 43372
rect 39228 43426 39284 43438
rect 39228 43374 39230 43426
rect 39282 43374 39284 43426
rect 39228 43316 39284 43374
rect 39228 43250 39284 43260
rect 39004 42756 39060 42766
rect 39452 42756 39508 42766
rect 39060 42754 39508 42756
rect 39060 42702 39454 42754
rect 39506 42702 39508 42754
rect 39060 42700 39508 42702
rect 39004 41970 39060 42700
rect 39452 42690 39508 42700
rect 39004 41918 39006 41970
rect 39058 41918 39060 41970
rect 39004 41906 39060 41918
rect 39228 42530 39284 42542
rect 39228 42478 39230 42530
rect 39282 42478 39284 42530
rect 39228 41748 39284 42478
rect 38780 41692 39284 41748
rect 39564 42532 39620 43596
rect 39900 42756 39956 42766
rect 39900 42662 39956 42700
rect 40012 42754 40068 42766
rect 40012 42702 40014 42754
rect 40066 42702 40068 42754
rect 40012 42532 40068 42702
rect 39564 42476 40068 42532
rect 40236 42754 40292 42766
rect 40236 42702 40238 42754
rect 40290 42702 40292 42754
rect 38444 40290 38500 40302
rect 38444 40238 38446 40290
rect 38498 40238 38500 40290
rect 38444 39844 38500 40238
rect 38444 39778 38500 39788
rect 38220 39730 38388 39732
rect 38220 39678 38222 39730
rect 38274 39678 38388 39730
rect 38220 39676 38388 39678
rect 38220 39666 38276 39676
rect 38332 39620 38388 39676
rect 38556 39620 38612 39630
rect 38332 39618 38612 39620
rect 38332 39566 38558 39618
rect 38610 39566 38612 39618
rect 38332 39564 38612 39566
rect 37996 39452 38276 39508
rect 37772 38274 37940 38276
rect 37772 38222 37774 38274
rect 37826 38222 37940 38274
rect 37772 38220 37940 38222
rect 37996 38612 38052 38622
rect 37772 38210 37828 38220
rect 36988 38108 37156 38164
rect 36988 37938 37044 37950
rect 36988 37886 36990 37938
rect 37042 37886 37044 37938
rect 36988 37604 37044 37886
rect 36988 37538 37044 37548
rect 36876 37326 36878 37378
rect 36930 37326 36932 37378
rect 36876 36932 36932 37326
rect 36988 37380 37044 37390
rect 37100 37380 37156 38108
rect 37884 37938 37940 37950
rect 37884 37886 37886 37938
rect 37938 37886 37940 37938
rect 37212 37828 37268 37838
rect 37212 37734 37268 37772
rect 37436 37828 37492 37838
rect 37884 37828 37940 37886
rect 37436 37826 37940 37828
rect 37436 37774 37438 37826
rect 37490 37774 37940 37826
rect 37436 37772 37940 37774
rect 37436 37762 37492 37772
rect 37212 37492 37268 37502
rect 37212 37490 37828 37492
rect 37212 37438 37214 37490
rect 37266 37438 37828 37490
rect 37212 37436 37828 37438
rect 37212 37426 37268 37436
rect 36988 37378 37156 37380
rect 36988 37326 36990 37378
rect 37042 37326 37156 37378
rect 36988 37324 37156 37326
rect 36988 37314 37044 37324
rect 36876 36866 36932 36876
rect 37100 36820 37156 37324
rect 37772 37154 37828 37436
rect 37772 37102 37774 37154
rect 37826 37102 37828 37154
rect 37772 37090 37828 37102
rect 37100 36764 37492 36820
rect 36876 36484 36932 36494
rect 36876 35922 36932 36428
rect 36876 35870 36878 35922
rect 36930 35870 36932 35922
rect 36876 35858 36932 35870
rect 36764 35196 37044 35252
rect 36036 35084 36372 35140
rect 35980 35074 36036 35084
rect 36316 35026 36372 35084
rect 36316 34974 36318 35026
rect 36370 34974 36372 35026
rect 36316 34962 36372 34974
rect 35868 34916 35924 34926
rect 35868 34822 35924 34860
rect 35532 34802 35700 34804
rect 35532 34750 35534 34802
rect 35586 34750 35700 34802
rect 35532 34748 35700 34750
rect 35532 34738 35588 34748
rect 36988 34132 37044 35196
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 33572 35252 33582
rect 35084 33570 35252 33572
rect 35084 33518 35198 33570
rect 35250 33518 35252 33570
rect 35084 33516 35252 33518
rect 35196 33506 35252 33516
rect 33068 33282 33124 33292
rect 35644 33348 35700 33358
rect 35644 33254 35700 33292
rect 36988 33346 37044 34076
rect 37324 34242 37380 34254
rect 37324 34190 37326 34242
rect 37378 34190 37380 34242
rect 37324 33348 37380 34190
rect 37436 33460 37492 36764
rect 37884 36708 37940 37772
rect 37996 37266 38052 38556
rect 37996 37214 37998 37266
rect 38050 37214 38052 37266
rect 37996 37202 38052 37214
rect 37884 36642 37940 36652
rect 37884 36484 37940 36494
rect 37884 36390 37940 36428
rect 37996 36372 38052 36382
rect 37996 36278 38052 36316
rect 37996 36148 38052 36158
rect 37772 33460 37828 33470
rect 37436 33458 37828 33460
rect 37436 33406 37438 33458
rect 37490 33406 37774 33458
rect 37826 33406 37828 33458
rect 37436 33404 37828 33406
rect 37436 33394 37492 33404
rect 37772 33394 37828 33404
rect 36988 33294 36990 33346
rect 37042 33294 37044 33346
rect 31836 33180 32004 33236
rect 31500 30930 31556 30940
rect 31612 32676 31668 32686
rect 30044 28642 30212 28644
rect 30044 28590 30046 28642
rect 30098 28590 30212 28642
rect 30044 28588 30212 28590
rect 30268 30210 30324 30222
rect 30268 30158 30270 30210
rect 30322 30158 30324 30210
rect 30268 28644 30324 30158
rect 31612 30100 31668 32620
rect 31836 32562 31892 33180
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32498 31892 32510
rect 34412 33122 34468 33134
rect 34412 33070 34414 33122
rect 34466 33070 34468 33122
rect 32956 30996 33012 31006
rect 33516 30996 33572 31006
rect 32956 30902 33012 30940
rect 33292 30994 33572 30996
rect 33292 30942 33518 30994
rect 33570 30942 33572 30994
rect 33292 30940 33572 30942
rect 31612 30034 31668 30044
rect 33068 30436 33124 30446
rect 32732 29986 32788 29998
rect 32732 29934 32734 29986
rect 32786 29934 32788 29986
rect 31276 29428 31332 29438
rect 30380 28644 30436 28654
rect 30324 28642 30436 28644
rect 30324 28590 30382 28642
rect 30434 28590 30436 28642
rect 30324 28588 30436 28590
rect 28476 27806 28478 27858
rect 28530 27806 28532 27858
rect 28476 27794 28532 27806
rect 30044 27858 30100 28588
rect 30268 28550 30324 28588
rect 30380 28578 30436 28588
rect 31276 28082 31332 29372
rect 32732 28532 32788 29934
rect 32732 28438 32788 28476
rect 31276 28030 31278 28082
rect 31330 28030 31332 28082
rect 31276 28018 31332 28030
rect 30940 27860 30996 27870
rect 30044 27806 30046 27858
rect 30098 27806 30100 27858
rect 30044 27794 30100 27806
rect 30828 27858 30996 27860
rect 30828 27806 30942 27858
rect 30994 27806 30996 27858
rect 30828 27804 30996 27806
rect 28140 27694 28142 27746
rect 28194 27694 28196 27746
rect 28140 27682 28196 27694
rect 30492 27748 30548 27758
rect 30828 27748 30884 27804
rect 30940 27794 30996 27804
rect 30492 27746 30884 27748
rect 30492 27694 30494 27746
rect 30546 27694 30884 27746
rect 30492 27692 30884 27694
rect 30492 27682 30548 27692
rect 27356 27634 27412 27646
rect 27356 27582 27358 27634
rect 27410 27582 27412 27634
rect 27356 27524 27412 27582
rect 26964 27468 27412 27524
rect 26908 27458 26964 27468
rect 26684 27134 26686 27186
rect 26738 27134 26740 27186
rect 26684 27122 26740 27134
rect 30828 26962 30884 27692
rect 30828 26910 30830 26962
rect 30882 26910 30884 26962
rect 30828 26908 30884 26910
rect 31724 27746 31780 27758
rect 31724 27694 31726 27746
rect 31778 27694 31780 27746
rect 30828 26852 30996 26908
rect 28364 26404 28420 26414
rect 30940 26404 30996 26852
rect 28364 26402 28532 26404
rect 28364 26350 28366 26402
rect 28418 26350 28532 26402
rect 28364 26348 28532 26350
rect 28364 26338 28420 26348
rect 26012 26126 26014 26178
rect 26066 26126 26068 26178
rect 26012 26114 26068 26126
rect 26124 26290 26180 26302
rect 28252 26292 28308 26302
rect 26124 26238 26126 26290
rect 26178 26238 26180 26290
rect 24780 25394 24836 25452
rect 25340 26068 25396 26078
rect 25340 25506 25396 26012
rect 26124 26068 26180 26238
rect 27916 26290 28308 26292
rect 27916 26238 28254 26290
rect 28306 26238 28308 26290
rect 27916 26236 28308 26238
rect 26124 26002 26180 26012
rect 26684 26180 26740 26190
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 25340 25442 25396 25454
rect 24780 25342 24782 25394
rect 24834 25342 24836 25394
rect 24780 25330 24836 25342
rect 25788 25396 25844 25406
rect 23660 24836 23716 24846
rect 23548 24834 23716 24836
rect 23548 24782 23662 24834
rect 23714 24782 23716 24834
rect 23548 24780 23716 24782
rect 23660 24770 23716 24780
rect 23324 24406 23380 24444
rect 23548 24500 23604 24510
rect 23548 24406 23604 24444
rect 22876 24098 22932 24108
rect 23324 24164 23380 24174
rect 21420 24052 21476 24062
rect 21420 23378 21476 23996
rect 22988 23940 23044 23950
rect 22988 23846 23044 23884
rect 22876 23828 22932 23838
rect 22876 23734 22932 23772
rect 21420 23326 21422 23378
rect 21474 23326 21476 23378
rect 21420 23156 21476 23326
rect 21420 23090 21476 23100
rect 21532 23714 21588 23726
rect 21532 23662 21534 23714
rect 21586 23662 21588 23714
rect 21532 22372 21588 23662
rect 21980 23714 22036 23726
rect 21980 23662 21982 23714
rect 22034 23662 22036 23714
rect 21980 23604 22036 23662
rect 21980 23538 22036 23548
rect 22652 23714 22708 23726
rect 23100 23716 23156 23726
rect 22652 23662 22654 23714
rect 22706 23662 22708 23714
rect 21980 23042 22036 23054
rect 21980 22990 21982 23042
rect 22034 22990 22036 23042
rect 21868 22930 21924 22942
rect 21868 22878 21870 22930
rect 21922 22878 21924 22930
rect 21532 22306 21588 22316
rect 21644 22372 21700 22382
rect 21644 22370 21812 22372
rect 21644 22318 21646 22370
rect 21698 22318 21812 22370
rect 21644 22316 21812 22318
rect 21644 22306 21700 22316
rect 21644 21812 21700 21822
rect 21644 21698 21700 21756
rect 21756 21810 21812 22316
rect 21756 21758 21758 21810
rect 21810 21758 21812 21810
rect 21756 21746 21812 21758
rect 21644 21646 21646 21698
rect 21698 21646 21700 21698
rect 21644 21634 21700 21646
rect 21868 21700 21924 22878
rect 21980 22484 22036 22990
rect 21980 22418 22036 22428
rect 22428 23042 22484 23054
rect 22428 22990 22430 23042
rect 22482 22990 22484 23042
rect 21980 22258 22036 22270
rect 21980 22206 21982 22258
rect 22034 22206 22036 22258
rect 21980 21810 22036 22206
rect 22428 21924 22484 22990
rect 22428 21858 22484 21868
rect 22540 23044 22596 23054
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 22316 21812 22372 21822
rect 21420 21474 21476 21486
rect 21420 21422 21422 21474
rect 21474 21422 21476 21474
rect 21084 20190 21086 20242
rect 21138 20190 21140 20242
rect 21084 20178 21140 20190
rect 21308 20690 21364 20702
rect 21308 20638 21310 20690
rect 21362 20638 21364 20690
rect 21308 20132 21364 20638
rect 21420 20468 21476 21422
rect 21868 20916 21924 21644
rect 22204 21698 22260 21710
rect 22204 21646 22206 21698
rect 22258 21646 22260 21698
rect 22204 21028 22260 21646
rect 22316 21698 22372 21756
rect 22316 21646 22318 21698
rect 22370 21646 22372 21698
rect 22316 21634 22372 21646
rect 22428 21028 22484 21038
rect 22204 20972 22428 21028
rect 22428 20962 22484 20972
rect 21868 20860 22260 20916
rect 21532 20692 21588 20702
rect 21532 20598 21588 20636
rect 21868 20690 21924 20702
rect 21868 20638 21870 20690
rect 21922 20638 21924 20690
rect 21420 20402 21476 20412
rect 21756 20578 21812 20590
rect 21756 20526 21758 20578
rect 21810 20526 21812 20578
rect 21756 20356 21812 20526
rect 21756 20290 21812 20300
rect 21308 20066 21364 20076
rect 21196 20018 21252 20030
rect 21196 19966 21198 20018
rect 21250 19966 21252 20018
rect 21196 18562 21252 19966
rect 21532 20020 21588 20030
rect 21532 19926 21588 19964
rect 21868 19908 21924 20638
rect 22092 20580 22148 20590
rect 21644 19852 21924 19908
rect 21980 20578 22148 20580
rect 21980 20526 22094 20578
rect 22146 20526 22148 20578
rect 21980 20524 22148 20526
rect 21308 19684 21364 19694
rect 21308 19458 21364 19628
rect 21308 19406 21310 19458
rect 21362 19406 21364 19458
rect 21308 19394 21364 19406
rect 21644 19458 21700 19852
rect 21644 19406 21646 19458
rect 21698 19406 21700 19458
rect 21644 19394 21700 19406
rect 21532 19348 21588 19358
rect 21532 19122 21588 19292
rect 21980 19346 22036 20524
rect 22092 20514 22148 20524
rect 21980 19294 21982 19346
rect 22034 19294 22036 19346
rect 21980 19282 22036 19294
rect 22092 19572 22148 19582
rect 21532 19070 21534 19122
rect 21586 19070 21588 19122
rect 21532 19058 21588 19070
rect 21756 19012 21812 19022
rect 21196 18510 21198 18562
rect 21250 18510 21252 18562
rect 21196 18498 21252 18510
rect 21308 18564 21364 18574
rect 21308 17444 21364 18508
rect 21756 18450 21812 18956
rect 21756 18398 21758 18450
rect 21810 18398 21812 18450
rect 21756 18386 21812 18398
rect 21980 18452 22036 18462
rect 21756 18228 21812 18238
rect 21532 18004 21588 18014
rect 21588 17948 21700 18004
rect 21532 17938 21588 17948
rect 21420 17668 21476 17678
rect 21420 17666 21588 17668
rect 21420 17614 21422 17666
rect 21474 17614 21588 17666
rect 21420 17612 21588 17614
rect 21420 17602 21476 17612
rect 21308 17388 21476 17444
rect 20860 16370 20916 16380
rect 21196 17220 21252 17230
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 20524 16034 20580 16046
rect 20972 16324 21028 16334
rect 20412 15374 20414 15426
rect 20466 15374 20468 15426
rect 20412 15362 20468 15374
rect 20188 14802 20244 14812
rect 20524 15314 20580 15326
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 19852 14690 19908 14700
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 14466 19796 14478
rect 19852 14418 19908 14430
rect 19852 14366 19854 14418
rect 19906 14366 19908 14418
rect 19740 14308 19796 14318
rect 19852 14308 19908 14366
rect 19796 14252 19908 14308
rect 20188 14306 20244 14318
rect 20188 14254 20190 14306
rect 20242 14254 20244 14306
rect 19740 14242 19796 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13916 19796 13972
rect 19516 13746 19572 13758
rect 19516 13694 19518 13746
rect 19570 13694 19572 13746
rect 19292 11442 19348 11452
rect 19404 13636 19460 13646
rect 19180 11342 19182 11394
rect 19234 11342 19236 11394
rect 19180 11330 19236 11342
rect 19068 10948 19124 10958
rect 19068 10276 19124 10892
rect 19180 10724 19236 10734
rect 19180 10610 19236 10668
rect 19180 10558 19182 10610
rect 19234 10558 19236 10610
rect 19180 10546 19236 10558
rect 19292 10612 19348 10622
rect 19068 10210 19124 10220
rect 19068 9156 19124 9166
rect 19068 8370 19124 9100
rect 19068 8318 19070 8370
rect 19122 8318 19124 8370
rect 19068 8306 19124 8318
rect 19292 8482 19348 10556
rect 19404 10386 19460 13580
rect 19516 12068 19572 13694
rect 19740 12850 19796 13916
rect 19852 13860 19908 13870
rect 19852 13076 19908 13804
rect 19852 12962 19908 13020
rect 19852 12910 19854 12962
rect 19906 12910 19908 12962
rect 19852 12898 19908 12910
rect 19740 12798 19742 12850
rect 19794 12798 19796 12850
rect 19740 12786 19796 12798
rect 20188 12740 20244 14254
rect 20524 14196 20580 15262
rect 20972 15148 21028 16268
rect 21196 15148 21252 17164
rect 21308 15876 21364 15886
rect 21308 15782 21364 15820
rect 21420 15316 21476 17388
rect 21532 16436 21588 17612
rect 21644 17554 21700 17948
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21644 17490 21700 17502
rect 21756 17220 21812 18172
rect 21980 17554 22036 18396
rect 22092 18116 22148 19516
rect 22204 18900 22260 20860
rect 22540 20804 22596 22988
rect 22652 21586 22708 23662
rect 22988 23660 23100 23716
rect 22988 23604 23044 23660
rect 23100 23622 23156 23660
rect 22876 23548 23044 23604
rect 22764 23154 22820 23166
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 22764 23042 22820 23102
rect 22764 22990 22766 23042
rect 22818 22990 22820 23042
rect 22764 22978 22820 22990
rect 22764 21812 22820 21822
rect 22876 21812 22932 23548
rect 23324 23492 23380 24108
rect 23548 23940 23604 23950
rect 23548 23938 23716 23940
rect 23548 23886 23550 23938
rect 23602 23886 23716 23938
rect 23548 23884 23716 23886
rect 23548 23874 23604 23884
rect 23660 23604 23716 23884
rect 23772 23828 23828 23838
rect 23884 23828 23940 25116
rect 25004 25282 25060 25294
rect 25004 25230 25006 25282
rect 25058 25230 25060 25282
rect 25004 24724 25060 25230
rect 25788 24946 25844 25340
rect 25788 24894 25790 24946
rect 25842 24894 25844 24946
rect 25788 24882 25844 24894
rect 25004 24658 25060 24668
rect 26012 24724 26068 24734
rect 25340 24612 25396 24622
rect 25676 24612 25732 24622
rect 25340 24610 25732 24612
rect 25340 24558 25342 24610
rect 25394 24558 25678 24610
rect 25730 24558 25732 24610
rect 25340 24556 25732 24558
rect 26012 24612 26068 24668
rect 26460 24612 26516 24622
rect 26012 24610 26628 24612
rect 26012 24558 26462 24610
rect 26514 24558 26628 24610
rect 26012 24556 26628 24558
rect 24556 24500 24612 24510
rect 24612 24444 24724 24500
rect 24556 24434 24612 24444
rect 23828 23772 23940 23828
rect 23772 23734 23828 23772
rect 24332 23714 24388 23726
rect 24332 23662 24334 23714
rect 24386 23662 24388 23714
rect 24332 23604 24388 23662
rect 23660 23548 24388 23604
rect 23660 23492 23716 23548
rect 23324 23436 23492 23492
rect 22820 21810 22932 21812
rect 22820 21758 22878 21810
rect 22930 21758 22932 21810
rect 22820 21756 22932 21758
rect 22764 21746 22820 21756
rect 22876 21746 22932 21756
rect 22988 21812 23044 21822
rect 22988 21718 23044 21756
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 21252 22708 21534
rect 23100 21588 23156 21598
rect 23100 21586 23268 21588
rect 23100 21534 23102 21586
rect 23154 21534 23268 21586
rect 23100 21532 23268 21534
rect 23100 21522 23156 21532
rect 22652 21186 22708 21196
rect 23100 21252 23156 21262
rect 22876 21028 22932 21038
rect 22876 20914 22932 20972
rect 22876 20862 22878 20914
rect 22930 20862 22932 20914
rect 22876 20850 22932 20862
rect 22540 20748 22820 20804
rect 22428 20690 22484 20702
rect 22428 20638 22430 20690
rect 22482 20638 22484 20690
rect 22316 20578 22372 20590
rect 22316 20526 22318 20578
rect 22370 20526 22372 20578
rect 22316 20468 22372 20526
rect 22316 19012 22372 20412
rect 22428 19572 22484 20638
rect 22764 19572 22820 20748
rect 23100 20020 23156 21196
rect 23212 20244 23268 21532
rect 23324 21586 23380 21598
rect 23324 21534 23326 21586
rect 23378 21534 23380 21586
rect 23324 20578 23380 21534
rect 23324 20526 23326 20578
rect 23378 20526 23380 20578
rect 23324 20468 23380 20526
rect 23324 20402 23380 20412
rect 23212 20178 23268 20188
rect 23324 20020 23380 20030
rect 23100 20018 23380 20020
rect 23100 19966 23326 20018
rect 23378 19966 23380 20018
rect 23100 19964 23380 19966
rect 23324 19954 23380 19964
rect 22428 19516 22708 19572
rect 22428 19348 22484 19358
rect 22428 19234 22484 19292
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 22428 19170 22484 19182
rect 22316 18956 22596 19012
rect 22204 18844 22484 18900
rect 22092 18060 22260 18116
rect 21980 17502 21982 17554
rect 22034 17502 22036 17554
rect 21980 17490 22036 17502
rect 21868 17444 21924 17454
rect 21868 17332 21924 17388
rect 21868 17276 22036 17332
rect 21756 17164 21924 17220
rect 21532 16380 21812 16436
rect 21644 16210 21700 16222
rect 21644 16158 21646 16210
rect 21698 16158 21700 16210
rect 21420 15222 21476 15260
rect 21532 15874 21588 15886
rect 21532 15822 21534 15874
rect 21586 15822 21588 15874
rect 20972 15092 21140 15148
rect 21196 15092 21476 15148
rect 20524 14140 20692 14196
rect 20524 13746 20580 13758
rect 20524 13694 20526 13746
rect 20578 13694 20580 13746
rect 20412 13524 20468 13534
rect 20188 12674 20244 12684
rect 20300 13522 20468 13524
rect 20300 13470 20414 13522
rect 20466 13470 20468 13522
rect 20300 13468 20468 13470
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19852 12292 19908 12302
rect 19852 12178 19908 12236
rect 19852 12126 19854 12178
rect 19906 12126 19908 12178
rect 19740 12068 19796 12078
rect 19516 12066 19796 12068
rect 19516 12014 19742 12066
rect 19794 12014 19796 12066
rect 19516 12012 19796 12014
rect 19740 12002 19796 12012
rect 19852 11788 19908 12126
rect 19628 11732 19908 11788
rect 20076 11844 20132 11854
rect 19628 10388 19684 11732
rect 20076 11618 20132 11788
rect 20076 11566 20078 11618
rect 20130 11566 20132 11618
rect 20076 11554 20132 11566
rect 19852 11508 19908 11518
rect 19908 11452 20020 11508
rect 19852 11442 19908 11452
rect 19964 11394 20020 11452
rect 19964 11342 19966 11394
rect 20018 11342 20020 11394
rect 19964 11330 20020 11342
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19404 10334 19406 10386
rect 19458 10334 19460 10386
rect 19404 10322 19460 10334
rect 19516 10332 19684 10388
rect 19740 10610 19796 10622
rect 19740 10558 19742 10610
rect 19794 10558 19796 10610
rect 19740 10388 19796 10558
rect 19516 9042 19572 10332
rect 19740 10322 19796 10332
rect 20188 10500 20244 10510
rect 20188 9938 20244 10444
rect 20188 9886 20190 9938
rect 20242 9886 20244 9938
rect 20188 9874 20244 9886
rect 19516 8990 19518 9042
rect 19570 8990 19572 9042
rect 19516 8978 19572 8990
rect 19628 9826 19684 9838
rect 19628 9774 19630 9826
rect 19682 9774 19684 9826
rect 19628 8932 19684 9774
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 8876 20020 8932
rect 19516 8820 19572 8830
rect 19516 8726 19572 8764
rect 19292 8430 19294 8482
rect 19346 8430 19348 8482
rect 18732 8206 18734 8258
rect 18786 8206 18788 8258
rect 18732 8194 18788 8206
rect 18844 8260 18900 8270
rect 17948 7646 17950 7698
rect 18002 7646 18004 7698
rect 17948 7634 18004 7646
rect 18060 8092 18340 8148
rect 17836 7586 17892 7598
rect 17836 7534 17838 7586
rect 17890 7534 17892 7586
rect 17836 7364 17892 7534
rect 17836 7298 17892 7308
rect 18060 6020 18116 8092
rect 18508 7364 18564 7374
rect 18508 7270 18564 7308
rect 18732 7252 18788 7262
rect 18396 6692 18452 6702
rect 18060 5926 18116 5964
rect 18284 6580 18340 6590
rect 17836 5908 17892 5918
rect 17836 5906 18004 5908
rect 17836 5854 17838 5906
rect 17890 5854 18004 5906
rect 17836 5852 18004 5854
rect 17836 5842 17892 5852
rect 17724 5628 17892 5684
rect 17724 4564 17780 4574
rect 17724 4470 17780 4508
rect 17612 4398 17614 4450
rect 17666 4398 17668 4450
rect 17612 4386 17668 4398
rect 17724 3668 17780 3678
rect 17724 3574 17780 3612
rect 17500 3332 17780 3388
rect 17276 3042 17332 3052
rect 15932 2930 15988 2940
rect 15372 2884 15428 2894
rect 15260 2828 15372 2884
rect 15372 2818 15428 2828
rect 15148 2706 15204 2716
rect 17724 2660 17780 3332
rect 17836 3220 17892 5628
rect 17948 5460 18004 5852
rect 17948 5124 18004 5404
rect 18284 5348 18340 6524
rect 18396 5684 18452 6636
rect 18396 5618 18452 5628
rect 18620 5572 18676 5582
rect 18284 5292 18564 5348
rect 18284 5124 18340 5134
rect 17948 5068 18284 5124
rect 18284 5030 18340 5068
rect 18060 4900 18116 4910
rect 18060 4806 18116 4844
rect 18172 4898 18228 4910
rect 18172 4846 18174 4898
rect 18226 4846 18228 4898
rect 18172 4564 18228 4846
rect 17948 4508 18228 4564
rect 18284 4788 18340 4798
rect 17948 4450 18004 4508
rect 17948 4398 17950 4450
rect 18002 4398 18004 4450
rect 17948 4386 18004 4398
rect 17836 3154 17892 3164
rect 18060 4340 18116 4350
rect 18284 4340 18340 4732
rect 18060 4338 18340 4340
rect 18060 4286 18062 4338
rect 18114 4286 18340 4338
rect 18060 4284 18340 4286
rect 17724 2594 17780 2604
rect 18060 2548 18116 4284
rect 18396 3668 18452 5292
rect 18508 5010 18564 5292
rect 18508 4958 18510 5010
rect 18562 4958 18564 5010
rect 18508 4946 18564 4958
rect 18396 3602 18452 3612
rect 18508 4564 18564 4574
rect 18620 4564 18676 5516
rect 18564 4508 18676 4564
rect 18508 3666 18564 4508
rect 18508 3614 18510 3666
rect 18562 3614 18564 3666
rect 18508 3602 18564 3614
rect 18732 3388 18788 7196
rect 18844 6132 18900 8204
rect 19292 8260 19348 8430
rect 19964 8482 20020 8876
rect 19964 8430 19966 8482
rect 20018 8430 20020 8482
rect 19964 8418 20020 8430
rect 20300 8428 20356 13468
rect 20412 13458 20468 13468
rect 20524 13076 20580 13694
rect 20412 13020 20580 13076
rect 20412 11844 20468 13020
rect 20636 12964 20692 14140
rect 20636 12870 20692 12908
rect 20972 13746 21028 13758
rect 20972 13694 20974 13746
rect 21026 13694 21028 13746
rect 20636 12740 20692 12750
rect 20972 12740 21028 13694
rect 20636 12738 21028 12740
rect 20636 12686 20638 12738
rect 20690 12686 21028 12738
rect 20636 12684 21028 12686
rect 20636 12674 20692 12684
rect 20412 11778 20468 11788
rect 20524 12628 20580 12638
rect 20524 10836 20580 12572
rect 20748 12180 20804 12190
rect 21084 12180 21140 15092
rect 21308 14756 21364 14766
rect 21196 14700 21308 14756
rect 21196 14530 21252 14700
rect 21308 14690 21364 14700
rect 21196 14478 21198 14530
rect 21250 14478 21252 14530
rect 21196 14466 21252 14478
rect 21420 14418 21476 15092
rect 21532 14868 21588 15822
rect 21532 14802 21588 14812
rect 21532 14532 21588 14542
rect 21644 14532 21700 16158
rect 21756 16098 21812 16380
rect 21756 16046 21758 16098
rect 21810 16046 21812 16098
rect 21756 15426 21812 16046
rect 21756 15374 21758 15426
rect 21810 15374 21812 15426
rect 21756 15362 21812 15374
rect 21532 14530 21700 14532
rect 21532 14478 21534 14530
rect 21586 14478 21700 14530
rect 21532 14476 21700 14478
rect 21756 15202 21812 15214
rect 21756 15150 21758 15202
rect 21810 15150 21812 15202
rect 21532 14466 21588 14476
rect 21420 14366 21422 14418
rect 21474 14366 21476 14418
rect 21420 14354 21476 14366
rect 21196 13636 21252 13646
rect 21196 13542 21252 13580
rect 21756 13524 21812 15150
rect 21532 13468 21812 13524
rect 21868 14418 21924 17164
rect 21868 14366 21870 14418
rect 21922 14366 21924 14418
rect 21196 13076 21252 13086
rect 21196 12516 21252 13020
rect 21420 12962 21476 12974
rect 21420 12910 21422 12962
rect 21474 12910 21476 12962
rect 21196 12460 21364 12516
rect 21196 12180 21252 12190
rect 21084 12178 21252 12180
rect 21084 12126 21198 12178
rect 21250 12126 21252 12178
rect 21084 12124 21252 12126
rect 20748 12086 20804 12124
rect 21196 12114 21252 12124
rect 20524 10770 20580 10780
rect 20636 11844 20692 11854
rect 20412 10612 20468 10622
rect 20412 10050 20468 10556
rect 20412 9998 20414 10050
rect 20466 9998 20468 10050
rect 20412 9986 20468 9998
rect 20524 10052 20580 10062
rect 20412 9828 20468 9838
rect 20524 9828 20580 9996
rect 20412 9826 20580 9828
rect 20412 9774 20414 9826
rect 20466 9774 20580 9826
rect 20412 9772 20580 9774
rect 20412 8596 20468 9772
rect 20636 9156 20692 11788
rect 21308 11394 21364 12460
rect 21420 12292 21476 12910
rect 21420 12226 21476 12236
rect 21308 11342 21310 11394
rect 21362 11342 21364 11394
rect 21308 11330 21364 11342
rect 20748 11170 20804 11182
rect 20748 11118 20750 11170
rect 20802 11118 20804 11170
rect 20748 10948 20804 11118
rect 20748 10882 20804 10892
rect 20860 10722 20916 10734
rect 20860 10670 20862 10722
rect 20914 10670 20916 10722
rect 20860 9940 20916 10670
rect 20860 9874 20916 9884
rect 20972 10610 21028 10622
rect 20972 10558 20974 10610
rect 21026 10558 21028 10610
rect 20748 9156 20804 9166
rect 20636 9154 20804 9156
rect 20636 9102 20750 9154
rect 20802 9102 20804 9154
rect 20636 9100 20804 9102
rect 20748 9090 20804 9100
rect 20524 8930 20580 8942
rect 20524 8878 20526 8930
rect 20578 8878 20580 8930
rect 20524 8708 20580 8878
rect 20524 8642 20580 8652
rect 20412 8530 20468 8540
rect 20300 8372 20468 8428
rect 19292 8194 19348 8204
rect 19516 8258 19572 8270
rect 19516 8206 19518 8258
rect 19570 8206 19572 8258
rect 19516 8036 19572 8206
rect 20188 8148 20244 8158
rect 20188 8054 20244 8092
rect 19516 7970 19572 7980
rect 19068 7924 19124 7934
rect 20300 7924 20356 7934
rect 19068 7700 19124 7868
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19068 7698 19348 7700
rect 19068 7646 19070 7698
rect 19122 7646 19348 7698
rect 19068 7644 19348 7646
rect 19068 7634 19124 7644
rect 19180 7252 19236 7262
rect 18956 7140 19012 7150
rect 18956 6690 19012 7084
rect 18956 6638 18958 6690
rect 19010 6638 19012 6690
rect 18956 6356 19012 6638
rect 18956 6290 19012 6300
rect 19180 7028 19236 7196
rect 19180 6244 19236 6972
rect 19292 6690 19348 7644
rect 20300 7698 20356 7868
rect 20300 7646 20302 7698
rect 20354 7646 20356 7698
rect 20300 7634 20356 7646
rect 20300 7476 20356 7486
rect 19740 7362 19796 7374
rect 19740 7310 19742 7362
rect 19794 7310 19796 7362
rect 19740 7252 19796 7310
rect 19740 7196 20020 7252
rect 19292 6638 19294 6690
rect 19346 6638 19348 6690
rect 19292 6626 19348 6638
rect 19852 6916 19908 6926
rect 19852 6690 19908 6860
rect 19852 6638 19854 6690
rect 19906 6638 19908 6690
rect 19852 6626 19908 6638
rect 19964 6692 20020 7196
rect 20188 7028 20244 7038
rect 19964 6626 20020 6636
rect 20076 6972 20188 7028
rect 20076 6578 20132 6972
rect 20188 6962 20244 6972
rect 20076 6526 20078 6578
rect 20130 6526 20132 6578
rect 20076 6514 20132 6526
rect 20188 6802 20244 6814
rect 20188 6750 20190 6802
rect 20242 6750 20244 6802
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19180 6188 19348 6244
rect 19836 6234 20100 6244
rect 18844 6076 19012 6132
rect 18844 5794 18900 5806
rect 18844 5742 18846 5794
rect 18898 5742 18900 5794
rect 18844 5684 18900 5742
rect 18844 5618 18900 5628
rect 18956 5460 19012 6076
rect 19180 6020 19236 6030
rect 19068 5906 19124 5918
rect 19068 5854 19070 5906
rect 19122 5854 19124 5906
rect 19068 5796 19124 5854
rect 19068 5730 19124 5740
rect 18844 5404 19012 5460
rect 19068 5572 19124 5582
rect 18844 4450 18900 5404
rect 19068 5122 19124 5516
rect 19068 5070 19070 5122
rect 19122 5070 19124 5122
rect 19068 5058 19124 5070
rect 19180 4788 19236 5964
rect 19292 5908 19348 6188
rect 19404 6132 19460 6142
rect 19404 6038 19460 6076
rect 19292 5852 19460 5908
rect 18844 4398 18846 4450
rect 18898 4398 18900 4450
rect 18844 4386 18900 4398
rect 19068 4732 19236 4788
rect 19292 4900 19348 4910
rect 18956 4228 19012 4238
rect 18956 4134 19012 4172
rect 18956 3668 19012 3678
rect 18732 3332 18900 3388
rect 18060 2482 18116 2492
rect 14924 2146 14980 2156
rect 18844 1652 18900 3332
rect 18956 2772 19012 3612
rect 19068 3332 19124 4732
rect 19292 4340 19348 4844
rect 19292 4246 19348 4284
rect 19180 4114 19236 4126
rect 19180 4062 19182 4114
rect 19234 4062 19236 4114
rect 19180 4004 19236 4062
rect 19180 3556 19236 3948
rect 19404 3666 19460 5852
rect 20188 5906 20244 6750
rect 20188 5854 20190 5906
rect 20242 5854 20244 5906
rect 20188 5842 20244 5854
rect 19740 5796 19796 5806
rect 19628 5794 19796 5796
rect 19628 5742 19742 5794
rect 19794 5742 19796 5794
rect 19628 5740 19796 5742
rect 19628 5348 19684 5740
rect 19740 5730 19796 5740
rect 19516 4788 19572 4798
rect 19628 4788 19684 5292
rect 20300 5122 20356 7420
rect 20412 6132 20468 8372
rect 20636 8370 20692 8382
rect 20636 8318 20638 8370
rect 20690 8318 20692 8370
rect 20524 7588 20580 7598
rect 20524 7494 20580 7532
rect 20636 7586 20692 8318
rect 20636 7534 20638 7586
rect 20690 7534 20692 7586
rect 20636 7476 20692 7534
rect 20636 7410 20692 7420
rect 20636 7250 20692 7262
rect 20636 7198 20638 7250
rect 20690 7198 20692 7250
rect 20412 6076 20580 6132
rect 20300 5070 20302 5122
rect 20354 5070 20356 5122
rect 20300 5058 20356 5070
rect 20412 5572 20468 5582
rect 19572 4732 19684 4788
rect 19836 4732 20100 4742
rect 19516 4722 19572 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19964 4340 20020 4350
rect 19964 4246 20020 4284
rect 19404 3614 19406 3666
rect 19458 3614 19460 3666
rect 19404 3602 19460 3614
rect 20300 3780 20356 3790
rect 20412 3780 20468 5516
rect 20356 3724 20468 3780
rect 20300 3666 20356 3724
rect 20300 3614 20302 3666
rect 20354 3614 20356 3666
rect 20300 3602 20356 3614
rect 19180 3490 19236 3500
rect 19852 3444 19908 3482
rect 20524 3388 20580 6076
rect 20636 5908 20692 7198
rect 20636 5842 20692 5852
rect 20860 5684 20916 5694
rect 20972 5684 21028 10558
rect 21308 10276 21364 10286
rect 21084 9828 21140 9838
rect 21084 9042 21140 9772
rect 21084 8990 21086 9042
rect 21138 8990 21140 9042
rect 21084 8484 21140 8990
rect 21084 8418 21140 8428
rect 21196 9492 21252 9502
rect 21084 8148 21140 8158
rect 21084 7252 21140 8092
rect 21084 7186 21140 7196
rect 21196 7028 21252 9436
rect 21308 7588 21364 10220
rect 21532 9044 21588 13468
rect 21868 13300 21924 14366
rect 21644 13244 21924 13300
rect 21644 11788 21700 13244
rect 21868 12964 21924 12974
rect 21868 12870 21924 12908
rect 21980 11956 22036 17276
rect 22204 16772 22260 18060
rect 22204 16706 22260 16716
rect 22428 16770 22484 18844
rect 22540 18228 22596 18956
rect 22540 18162 22596 18172
rect 22540 17554 22596 17566
rect 22540 17502 22542 17554
rect 22594 17502 22596 17554
rect 22540 17108 22596 17502
rect 22540 17042 22596 17052
rect 22428 16718 22430 16770
rect 22482 16718 22484 16770
rect 22092 15988 22148 15998
rect 22092 15894 22148 15932
rect 22316 15876 22372 15886
rect 22204 15820 22316 15876
rect 22204 15428 22260 15820
rect 22316 15810 22372 15820
rect 22092 15372 22260 15428
rect 22316 15652 22372 15662
rect 22092 12180 22148 15372
rect 22316 14530 22372 15596
rect 22316 14478 22318 14530
rect 22370 14478 22372 14530
rect 22316 14466 22372 14478
rect 22316 12852 22372 12862
rect 22092 12114 22148 12124
rect 22204 12850 22372 12852
rect 22204 12798 22318 12850
rect 22370 12798 22372 12850
rect 22204 12796 22372 12798
rect 21980 11890 22036 11900
rect 21868 11844 21924 11854
rect 21644 11732 21812 11788
rect 21644 11508 21700 11518
rect 21644 10834 21700 11452
rect 21644 10782 21646 10834
rect 21698 10782 21700 10834
rect 21644 10770 21700 10782
rect 21756 10612 21812 11732
rect 21868 11506 21924 11788
rect 22204 11620 22260 12796
rect 22316 12786 22372 12796
rect 21868 11454 21870 11506
rect 21922 11454 21924 11506
rect 21868 11442 21924 11454
rect 21980 11564 22260 11620
rect 22316 12068 22372 12078
rect 21644 10556 21812 10612
rect 21644 9604 21700 10556
rect 21756 9828 21812 9838
rect 21756 9734 21812 9772
rect 21644 9548 21812 9604
rect 21532 8978 21588 8988
rect 21420 8930 21476 8942
rect 21420 8878 21422 8930
rect 21474 8878 21476 8930
rect 21420 8260 21476 8878
rect 21420 8194 21476 8204
rect 21644 8148 21700 8158
rect 21644 8054 21700 8092
rect 21308 7532 21700 7588
rect 20916 5628 21028 5684
rect 21084 6972 21252 7028
rect 21308 7362 21364 7374
rect 21308 7310 21310 7362
rect 21362 7310 21364 7362
rect 21308 7028 21364 7310
rect 20860 5122 20916 5628
rect 20860 5070 20862 5122
rect 20914 5070 20916 5122
rect 20860 4788 20916 5070
rect 20860 4722 20916 4732
rect 20972 4900 21028 4910
rect 21084 4900 21140 6972
rect 21308 6962 21364 6972
rect 21196 6804 21252 6814
rect 21196 5236 21252 6748
rect 21308 6692 21364 6702
rect 21308 5906 21364 6636
rect 21420 6690 21476 6702
rect 21420 6638 21422 6690
rect 21474 6638 21476 6690
rect 21420 6468 21476 6638
rect 21420 6402 21476 6412
rect 21532 6578 21588 6590
rect 21532 6526 21534 6578
rect 21586 6526 21588 6578
rect 21308 5854 21310 5906
rect 21362 5854 21364 5906
rect 21308 5460 21364 5854
rect 21308 5394 21364 5404
rect 21420 6244 21476 6254
rect 21420 5346 21476 6188
rect 21420 5294 21422 5346
rect 21474 5294 21476 5346
rect 21420 5282 21476 5294
rect 21532 5796 21588 6526
rect 21196 5170 21252 5180
rect 21308 5124 21364 5134
rect 21308 5030 21364 5068
rect 21420 5010 21476 5022
rect 21420 4958 21422 5010
rect 21474 4958 21476 5010
rect 21084 4844 21364 4900
rect 20972 4226 21028 4844
rect 20972 4174 20974 4226
rect 21026 4174 21028 4226
rect 20972 3892 21028 4174
rect 20972 3826 21028 3836
rect 21308 3666 21364 4844
rect 21420 4452 21476 4958
rect 21420 3892 21476 4396
rect 21532 4338 21588 5740
rect 21532 4286 21534 4338
rect 21586 4286 21588 4338
rect 21532 4274 21588 4286
rect 21420 3826 21476 3836
rect 21308 3614 21310 3666
rect 21362 3614 21364 3666
rect 21308 3602 21364 3614
rect 21644 3668 21700 7532
rect 21756 7362 21812 9548
rect 21868 9042 21924 9054
rect 21868 8990 21870 9042
rect 21922 8990 21924 9042
rect 21868 8932 21924 8990
rect 21868 8260 21924 8876
rect 21980 8484 22036 11564
rect 22204 10612 22260 10622
rect 22204 10518 22260 10556
rect 22204 10052 22260 10062
rect 22316 10052 22372 12012
rect 22428 11396 22484 16718
rect 22540 16772 22596 16782
rect 22540 15764 22596 16716
rect 22540 15426 22596 15708
rect 22652 16212 22708 19516
rect 22764 19506 22820 19516
rect 22764 19010 22820 19022
rect 23100 19012 23156 19022
rect 22764 18958 22766 19010
rect 22818 18958 22820 19010
rect 22764 16884 22820 18958
rect 22876 19010 23156 19012
rect 22876 18958 23102 19010
rect 23154 18958 23156 19010
rect 22876 18956 23156 18958
rect 22876 16996 22932 18956
rect 23100 18946 23156 18956
rect 23212 18452 23268 18462
rect 23100 18450 23268 18452
rect 23100 18398 23214 18450
rect 23266 18398 23268 18450
rect 23100 18396 23268 18398
rect 22988 17442 23044 17454
rect 22988 17390 22990 17442
rect 23042 17390 23044 17442
rect 22988 17332 23044 17390
rect 22988 17266 23044 17276
rect 22876 16940 23044 16996
rect 22764 16828 22932 16884
rect 22652 15652 22708 16156
rect 22764 16658 22820 16670
rect 22764 16606 22766 16658
rect 22818 16606 22820 16658
rect 22764 16100 22820 16606
rect 22764 16034 22820 16044
rect 22652 15586 22708 15596
rect 22540 15374 22542 15426
rect 22594 15374 22596 15426
rect 22540 15362 22596 15374
rect 22764 15316 22820 15354
rect 22764 15250 22820 15260
rect 22876 15148 22932 16828
rect 22988 16548 23044 16940
rect 22988 16482 23044 16492
rect 23100 15988 23156 18396
rect 23212 18386 23268 18396
rect 23436 18228 23492 23436
rect 23548 23436 23716 23492
rect 23548 21028 23604 23436
rect 24556 23380 24612 23390
rect 23884 23042 23940 23054
rect 23884 22990 23886 23042
rect 23938 22990 23940 23042
rect 23548 20962 23604 20972
rect 23660 22370 23716 22382
rect 23660 22318 23662 22370
rect 23714 22318 23716 22370
rect 23660 20132 23716 22318
rect 23772 21474 23828 21486
rect 23772 21422 23774 21474
rect 23826 21422 23828 21474
rect 23772 21252 23828 21422
rect 23772 21186 23828 21196
rect 23884 21140 23940 22990
rect 24332 22932 24388 22942
rect 23884 21074 23940 21084
rect 24108 21586 24164 21598
rect 24108 21534 24110 21586
rect 24162 21534 24164 21586
rect 23772 20916 23828 20926
rect 23772 20822 23828 20860
rect 24108 20916 24164 21534
rect 24332 21588 24388 22876
rect 24332 21494 24388 21532
rect 24444 22260 24500 22270
rect 24220 21476 24276 21486
rect 24220 21382 24276 21420
rect 24444 20916 24500 22204
rect 24556 21364 24612 23324
rect 24668 21924 24724 24444
rect 25340 24388 25396 24556
rect 25676 24546 25732 24556
rect 26460 24546 26516 24556
rect 25340 24322 25396 24332
rect 25228 24276 25284 24286
rect 25228 24050 25284 24220
rect 25228 23998 25230 24050
rect 25282 23998 25284 24050
rect 25004 23828 25060 23838
rect 25004 23734 25060 23772
rect 24892 23716 24948 23726
rect 24780 22372 24836 22382
rect 24780 22278 24836 22316
rect 24668 21858 24724 21868
rect 24556 21298 24612 21308
rect 24668 21588 24724 21598
rect 23772 20244 23828 20254
rect 24108 20244 24164 20860
rect 23828 20188 23940 20244
rect 23772 20178 23828 20188
rect 23660 19460 23716 20076
rect 23660 19394 23716 19404
rect 23772 19906 23828 19918
rect 23772 19854 23774 19906
rect 23826 19854 23828 19906
rect 23660 18900 23716 18910
rect 23212 18172 23492 18228
rect 23548 18844 23660 18900
rect 23212 17220 23268 18172
rect 23436 17556 23492 17594
rect 23548 17556 23604 18844
rect 23660 18834 23716 18844
rect 23660 18340 23716 18350
rect 23772 18340 23828 19854
rect 23660 18338 23828 18340
rect 23660 18286 23662 18338
rect 23714 18286 23828 18338
rect 23660 18284 23828 18286
rect 23660 17780 23716 18284
rect 23660 17714 23716 17724
rect 23772 17668 23828 17678
rect 23548 17500 23716 17556
rect 23436 17490 23492 17500
rect 23212 17164 23492 17220
rect 23212 16884 23268 16894
rect 23212 16790 23268 16828
rect 23436 16324 23492 17164
rect 23324 16268 23492 16324
rect 23548 16772 23604 16782
rect 23212 16100 23268 16110
rect 23212 16006 23268 16044
rect 23100 15428 23156 15932
rect 23100 15362 23156 15372
rect 22876 15092 23156 15148
rect 22988 14532 23044 14542
rect 22988 14438 23044 14476
rect 22764 14306 22820 14318
rect 22764 14254 22766 14306
rect 22818 14254 22820 14306
rect 22652 13412 22708 13422
rect 22540 13356 22652 13412
rect 22540 12850 22596 13356
rect 22652 13346 22708 13356
rect 22764 13300 22820 14254
rect 22764 13234 22820 13244
rect 22652 13076 22708 13086
rect 22652 13074 23044 13076
rect 22652 13022 22654 13074
rect 22706 13022 23044 13074
rect 22652 13020 23044 13022
rect 22652 13010 22708 13020
rect 22988 12962 23044 13020
rect 22988 12910 22990 12962
rect 23042 12910 23044 12962
rect 22988 12898 23044 12910
rect 22540 12798 22542 12850
rect 22594 12798 22596 12850
rect 22540 12786 22596 12798
rect 23100 12740 23156 15092
rect 23324 14532 23380 16268
rect 23436 15876 23492 15886
rect 23436 15538 23492 15820
rect 23436 15486 23438 15538
rect 23490 15486 23492 15538
rect 23436 15474 23492 15486
rect 23324 14466 23380 14476
rect 23436 14308 23492 14318
rect 23324 13746 23380 13758
rect 23324 13694 23326 13746
rect 23378 13694 23380 13746
rect 23324 13412 23380 13694
rect 22876 12684 23156 12740
rect 23212 13356 23324 13412
rect 22652 12292 22708 12302
rect 22428 11330 22484 11340
rect 22540 12180 22596 12190
rect 22540 10164 22596 12124
rect 22204 10050 22372 10052
rect 22204 9998 22206 10050
rect 22258 9998 22372 10050
rect 22204 9996 22372 9998
rect 22428 10108 22596 10164
rect 22092 9826 22148 9838
rect 22092 9774 22094 9826
rect 22146 9774 22148 9826
rect 22092 9156 22148 9774
rect 22204 9268 22260 9996
rect 22204 9202 22260 9212
rect 22092 9090 22148 9100
rect 21980 8418 22036 8428
rect 22092 8932 22148 8942
rect 21980 8260 22036 8270
rect 21868 8258 22036 8260
rect 21868 8206 21982 8258
rect 22034 8206 22036 8258
rect 21868 8204 22036 8206
rect 21980 8194 22036 8204
rect 22092 8036 22148 8876
rect 21756 7310 21758 7362
rect 21810 7310 21812 7362
rect 21756 6244 21812 7310
rect 21756 6178 21812 6188
rect 21868 7980 22148 8036
rect 22204 8820 22260 8830
rect 21868 4900 21924 7980
rect 22092 7476 22148 7486
rect 21980 7474 22148 7476
rect 21980 7422 22094 7474
rect 22146 7422 22148 7474
rect 21980 7420 22148 7422
rect 21980 5012 22036 7420
rect 22092 7410 22148 7420
rect 22092 6578 22148 6590
rect 22092 6526 22094 6578
rect 22146 6526 22148 6578
rect 22092 6020 22148 6526
rect 22092 5684 22148 5964
rect 22204 5906 22260 8764
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 22204 5842 22260 5854
rect 22316 8260 22372 8270
rect 22316 5796 22372 8204
rect 22428 6580 22484 10108
rect 22652 9826 22708 12236
rect 22764 12178 22820 12190
rect 22764 12126 22766 12178
rect 22818 12126 22820 12178
rect 22764 9940 22820 12126
rect 22764 9874 22820 9884
rect 22652 9774 22654 9826
rect 22706 9774 22708 9826
rect 22652 9762 22708 9774
rect 22876 9604 22932 12684
rect 23212 12068 23268 13356
rect 23324 13346 23380 13356
rect 23436 12964 23492 14252
rect 23436 12898 23492 12908
rect 23548 13746 23604 16716
rect 23660 15148 23716 17500
rect 23772 17332 23828 17612
rect 23772 17266 23828 17276
rect 23772 16996 23828 17006
rect 23884 16996 23940 20188
rect 24108 20178 24164 20188
rect 24332 20860 24500 20916
rect 24332 20130 24388 20860
rect 24556 20802 24612 20814
rect 24556 20750 24558 20802
rect 24610 20750 24612 20802
rect 24556 20356 24612 20750
rect 24668 20692 24724 21532
rect 24780 20692 24836 20702
rect 24668 20690 24836 20692
rect 24668 20638 24782 20690
rect 24834 20638 24836 20690
rect 24668 20636 24836 20638
rect 24780 20626 24836 20636
rect 24892 20580 24948 23660
rect 25228 22372 25284 23998
rect 26124 23940 26180 23950
rect 26012 23938 26180 23940
rect 26012 23886 26126 23938
rect 26178 23886 26180 23938
rect 26012 23884 26180 23886
rect 25564 23828 25620 23838
rect 25564 23734 25620 23772
rect 25340 23716 25396 23726
rect 25340 23622 25396 23660
rect 25676 23380 25732 23390
rect 25564 23268 25620 23278
rect 25676 23268 25732 23324
rect 25564 23266 25732 23268
rect 25564 23214 25566 23266
rect 25618 23214 25732 23266
rect 25564 23212 25732 23214
rect 25564 23202 25620 23212
rect 25676 23044 25732 23054
rect 26012 23044 26068 23884
rect 26124 23874 26180 23884
rect 26460 23828 26516 23838
rect 26124 23380 26180 23390
rect 26180 23324 26292 23380
rect 26124 23314 26180 23324
rect 25676 23042 26068 23044
rect 25676 22990 25678 23042
rect 25730 22990 26068 23042
rect 25676 22988 26068 22990
rect 26124 23044 26180 23054
rect 25676 22978 25732 22988
rect 26124 22950 26180 22988
rect 25340 22932 25396 22942
rect 25340 22838 25396 22876
rect 24556 20300 24836 20356
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24108 20018 24164 20030
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 23772 16994 23940 16996
rect 23772 16942 23774 16994
rect 23826 16942 23940 16994
rect 23772 16940 23940 16942
rect 23996 19906 24052 19918
rect 23996 19854 23998 19906
rect 24050 19854 24052 19906
rect 23772 16930 23828 16940
rect 23884 16772 23940 16782
rect 23884 16678 23940 16716
rect 23996 16436 24052 19854
rect 24108 19908 24164 19966
rect 24108 19842 24164 19852
rect 24332 19796 24388 20078
rect 24332 19730 24388 19740
rect 24780 19684 24836 20300
rect 24780 19618 24836 19628
rect 24332 19460 24388 19470
rect 24892 19460 24948 20524
rect 24332 19366 24388 19404
rect 24556 19404 24948 19460
rect 25004 22316 25284 22372
rect 24332 19012 24388 19022
rect 24332 18452 24388 18956
rect 24444 18676 24500 18686
rect 24444 18582 24500 18620
rect 24556 18674 24612 19404
rect 24892 19236 24948 19246
rect 25004 19236 25060 22316
rect 25452 22260 25508 22270
rect 25452 22166 25508 22204
rect 26124 22260 26180 22270
rect 26236 22260 26292 23324
rect 26124 22258 26292 22260
rect 26124 22206 26126 22258
rect 26178 22206 26292 22258
rect 26124 22204 26292 22206
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26124 22194 26180 22204
rect 25228 22148 25284 22158
rect 25228 22054 25284 22092
rect 25788 22146 25844 22158
rect 25788 22094 25790 22146
rect 25842 22094 25844 22146
rect 25116 21924 25172 21934
rect 25172 21868 25284 21924
rect 25116 21858 25172 21868
rect 24892 19234 25060 19236
rect 24892 19182 24894 19234
rect 24946 19182 25060 19234
rect 24892 19180 25060 19182
rect 25116 21252 25172 21262
rect 25116 20020 25172 21196
rect 24892 19170 24948 19180
rect 25116 19012 25172 19964
rect 24556 18622 24558 18674
rect 24610 18622 24612 18674
rect 24556 18610 24612 18622
rect 24892 18956 25172 19012
rect 25228 20804 25284 21868
rect 25340 21812 25396 21822
rect 25340 21718 25396 21756
rect 25340 21588 25396 21598
rect 25340 21252 25396 21532
rect 25788 21588 25844 22094
rect 26236 21700 26292 21710
rect 25788 21494 25844 21532
rect 26124 21586 26180 21598
rect 26124 21534 26126 21586
rect 26178 21534 26180 21586
rect 26124 21476 26180 21534
rect 26124 21410 26180 21420
rect 25900 21252 25956 21262
rect 25340 21196 25508 21252
rect 25340 20804 25396 20814
rect 25228 20802 25396 20804
rect 25228 20750 25342 20802
rect 25394 20750 25396 20802
rect 25228 20748 25396 20750
rect 24332 18396 24500 18452
rect 24332 18226 24388 18238
rect 24332 18174 24334 18226
rect 24386 18174 24388 18226
rect 24332 18116 24388 18174
rect 24108 18060 24388 18116
rect 24108 17892 24164 18060
rect 24332 17892 24388 17902
rect 24108 17836 24276 17892
rect 24108 17668 24164 17678
rect 24108 17554 24164 17612
rect 24108 17502 24110 17554
rect 24162 17502 24164 17554
rect 24108 17490 24164 17502
rect 24220 17556 24276 17836
rect 24108 16660 24164 16670
rect 24220 16660 24276 17500
rect 24164 16604 24276 16660
rect 24332 16882 24388 17836
rect 24444 17666 24500 18396
rect 24444 17614 24446 17666
rect 24498 17614 24500 17666
rect 24444 17602 24500 17614
rect 24780 17444 24836 17454
rect 24780 17350 24836 17388
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 24108 16566 24164 16604
rect 24332 16436 24388 16830
rect 23996 16380 24276 16436
rect 23660 15092 23828 15148
rect 23772 14642 23828 15092
rect 23772 14590 23774 14642
rect 23826 14590 23828 14642
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 23212 11974 23268 12012
rect 23324 12852 23380 12862
rect 23324 11954 23380 12796
rect 23324 11902 23326 11954
rect 23378 11902 23380 11954
rect 22988 11396 23044 11406
rect 22988 11282 23044 11340
rect 22988 11230 22990 11282
rect 23042 11230 23044 11282
rect 22988 10722 23044 11230
rect 22988 10670 22990 10722
rect 23042 10670 23044 10722
rect 22988 10658 23044 10670
rect 23100 9940 23156 9950
rect 23156 9884 23268 9940
rect 23100 9846 23156 9884
rect 22652 9548 22932 9604
rect 22988 9716 23044 9726
rect 22652 9266 22708 9548
rect 22652 9214 22654 9266
rect 22706 9214 22708 9266
rect 22652 9202 22708 9214
rect 22764 9268 22820 9278
rect 22764 9174 22820 9212
rect 22540 8820 22596 8830
rect 22764 8820 22820 8830
rect 22540 8818 22764 8820
rect 22540 8766 22542 8818
rect 22594 8766 22764 8818
rect 22540 8764 22764 8766
rect 22540 8754 22596 8764
rect 22764 8754 22820 8764
rect 22540 8258 22596 8270
rect 22540 8206 22542 8258
rect 22594 8206 22596 8258
rect 22540 8036 22596 8206
rect 22540 7970 22596 7980
rect 22652 7476 22708 7486
rect 22988 7476 23044 9660
rect 23100 8260 23156 8270
rect 23100 8166 23156 8204
rect 22652 7474 23044 7476
rect 22652 7422 22654 7474
rect 22706 7422 23044 7474
rect 22652 7420 23044 7422
rect 23212 7474 23268 9884
rect 23324 9380 23380 11902
rect 23548 11844 23604 13694
rect 23660 14418 23716 14430
rect 23660 14366 23662 14418
rect 23714 14366 23716 14418
rect 23660 11956 23716 14366
rect 23772 13972 23828 14590
rect 23772 13906 23828 13916
rect 23996 14530 24052 14542
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 23772 13634 23828 13646
rect 23772 13582 23774 13634
rect 23826 13582 23828 13634
rect 23772 12852 23828 13582
rect 23772 12786 23828 12796
rect 23884 13522 23940 13534
rect 23884 13470 23886 13522
rect 23938 13470 23940 13522
rect 23884 12180 23940 13470
rect 23884 12114 23940 12124
rect 23996 12962 24052 14478
rect 23996 12910 23998 12962
rect 24050 12910 24052 12962
rect 23660 11900 23940 11956
rect 23548 11788 23828 11844
rect 23436 11396 23492 11406
rect 23436 11394 23604 11396
rect 23436 11342 23438 11394
rect 23490 11342 23604 11394
rect 23436 11340 23604 11342
rect 23436 11330 23492 11340
rect 23324 9324 23492 9380
rect 23212 7422 23214 7474
rect 23266 7422 23268 7474
rect 22652 7410 22708 7420
rect 23212 7410 23268 7422
rect 23324 9156 23380 9166
rect 22540 6804 22596 6814
rect 22540 6710 22596 6748
rect 22988 6690 23044 6702
rect 22988 6638 22990 6690
rect 23042 6638 23044 6690
rect 22764 6580 22820 6590
rect 22428 6578 22932 6580
rect 22428 6526 22766 6578
rect 22818 6526 22932 6578
rect 22428 6524 22932 6526
rect 22764 6514 22820 6524
rect 22316 5740 22820 5796
rect 22092 5618 22148 5628
rect 22540 5236 22596 5246
rect 22540 5142 22596 5180
rect 22764 5122 22820 5740
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 21980 4956 22372 5012
rect 21868 4844 22260 4900
rect 21756 4338 21812 4350
rect 21756 4286 21758 4338
rect 21810 4286 21812 4338
rect 21756 4228 21812 4286
rect 21756 4162 21812 4172
rect 21756 3668 21812 3678
rect 21644 3666 21812 3668
rect 21644 3614 21758 3666
rect 21810 3614 21812 3666
rect 21644 3612 21812 3614
rect 21756 3602 21812 3612
rect 22092 3668 22148 3678
rect 22204 3668 22260 4844
rect 22316 4116 22372 4956
rect 22428 4116 22484 4126
rect 22316 4060 22428 4116
rect 22092 3666 22260 3668
rect 22092 3614 22094 3666
rect 22146 3614 22260 3666
rect 22092 3612 22260 3614
rect 22092 3602 22148 3612
rect 22428 3554 22484 4060
rect 22764 3668 22820 5070
rect 22764 3602 22820 3612
rect 22428 3502 22430 3554
rect 22482 3502 22484 3554
rect 22428 3490 22484 3502
rect 19068 3266 19124 3276
rect 19628 3332 19908 3388
rect 20412 3332 20580 3388
rect 22876 3332 22932 6524
rect 22988 6020 23044 6638
rect 22988 4114 23044 5964
rect 23100 5908 23156 5918
rect 23100 5814 23156 5852
rect 22988 4062 22990 4114
rect 23042 4062 23044 4114
rect 22988 4050 23044 4062
rect 23212 3444 23268 3482
rect 23324 3444 23380 9100
rect 23436 8820 23492 9324
rect 23436 8754 23492 8764
rect 23436 8036 23492 8046
rect 23436 7362 23492 7980
rect 23548 7586 23604 11340
rect 23660 9044 23716 9054
rect 23660 8950 23716 8988
rect 23660 8708 23716 8718
rect 23772 8708 23828 11788
rect 23884 11060 23940 11900
rect 23884 10612 23940 11004
rect 23884 10546 23940 10556
rect 23884 9826 23940 9838
rect 23884 9774 23886 9826
rect 23938 9774 23940 9826
rect 23884 9044 23940 9774
rect 23996 9268 24052 12910
rect 24108 13300 24164 13310
rect 24108 11956 24164 13244
rect 24220 12850 24276 16380
rect 24332 16370 24388 16380
rect 24780 17108 24836 17118
rect 24780 16212 24836 17052
rect 24556 16156 24836 16212
rect 24556 16098 24612 16156
rect 24556 16046 24558 16098
rect 24610 16046 24612 16098
rect 24556 16034 24612 16046
rect 24780 15988 24836 15998
rect 24332 15316 24388 15326
rect 24332 15222 24388 15260
rect 24556 15202 24612 15214
rect 24556 15150 24558 15202
rect 24610 15150 24612 15202
rect 24444 14530 24500 14542
rect 24444 14478 24446 14530
rect 24498 14478 24500 14530
rect 24444 14420 24500 14478
rect 24444 14354 24500 14364
rect 24220 12798 24222 12850
rect 24274 12798 24276 12850
rect 24220 12786 24276 12798
rect 24556 12852 24612 15150
rect 24668 15202 24724 15214
rect 24668 15150 24670 15202
rect 24722 15150 24724 15202
rect 24668 14644 24724 15150
rect 24668 14578 24724 14588
rect 24668 13972 24724 13982
rect 24780 13972 24836 15932
rect 24892 15148 24948 18956
rect 25116 17668 25172 17678
rect 25228 17668 25284 20748
rect 25340 20738 25396 20748
rect 25452 20690 25508 21196
rect 25452 20638 25454 20690
rect 25506 20638 25508 20690
rect 25452 20626 25508 20638
rect 25676 20692 25732 20702
rect 25676 20598 25732 20636
rect 25340 20020 25396 20030
rect 25676 20020 25732 20030
rect 25340 20018 25732 20020
rect 25340 19966 25342 20018
rect 25394 19966 25678 20018
rect 25730 19966 25732 20018
rect 25340 19964 25732 19966
rect 25340 19954 25396 19964
rect 25340 19572 25396 19582
rect 25396 19516 25508 19572
rect 25340 19506 25396 19516
rect 25340 19348 25396 19358
rect 25340 17892 25396 19292
rect 25452 18450 25508 19516
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 25452 18386 25508 18398
rect 25564 18452 25620 19964
rect 25676 19954 25732 19964
rect 25676 19796 25732 19806
rect 25676 18562 25732 19740
rect 25788 19234 25844 19246
rect 25788 19182 25790 19234
rect 25842 19182 25844 19234
rect 25788 19124 25844 19182
rect 25788 18676 25844 19068
rect 25900 18900 25956 21196
rect 25900 18834 25956 18844
rect 26124 20578 26180 20590
rect 26124 20526 26126 20578
rect 26178 20526 26180 20578
rect 26124 18676 26180 20526
rect 26236 20580 26292 21644
rect 26236 20514 26292 20524
rect 26236 20020 26292 20030
rect 26348 20020 26404 23102
rect 26460 20356 26516 23772
rect 26572 22372 26628 24556
rect 26684 23828 26740 26124
rect 26908 26178 26964 26190
rect 26908 26126 26910 26178
rect 26962 26126 26964 26178
rect 26908 26068 26964 26126
rect 27468 26180 27524 26190
rect 27468 26086 27524 26124
rect 26908 26002 26964 26012
rect 27244 26068 27300 26078
rect 27244 25284 27300 26012
rect 27916 25732 27972 26236
rect 28252 26226 28308 26236
rect 28364 26068 28420 26078
rect 28364 25974 28420 26012
rect 27916 25506 27972 25676
rect 27916 25454 27918 25506
rect 27970 25454 27972 25506
rect 27916 25442 27972 25454
rect 28252 25508 28308 25518
rect 28476 25508 28532 26348
rect 30940 26338 30996 26348
rect 31724 26404 31780 27694
rect 33068 27524 33124 30380
rect 33292 30210 33348 30940
rect 33516 30930 33572 30940
rect 33292 30158 33294 30210
rect 33346 30158 33348 30210
rect 33292 30146 33348 30158
rect 34300 30212 34356 30222
rect 33404 29538 33460 29550
rect 33404 29486 33406 29538
rect 33458 29486 33460 29538
rect 33180 27858 33236 27870
rect 33180 27806 33182 27858
rect 33234 27806 33236 27858
rect 33180 27748 33236 27806
rect 33180 27682 33236 27692
rect 33404 27860 33460 29486
rect 33628 29428 33684 29438
rect 33628 29334 33684 29372
rect 34300 28754 34356 30156
rect 34300 28702 34302 28754
rect 34354 28702 34356 28754
rect 34300 28690 34356 28702
rect 34412 29652 34468 33070
rect 36876 32676 36932 32686
rect 36876 32582 36932 32620
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35868 31108 35924 31118
rect 35756 31106 35924 31108
rect 35756 31054 35870 31106
rect 35922 31054 35924 31106
rect 35756 31052 35924 31054
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34748 30212 34804 30222
rect 34748 30118 34804 30156
rect 35532 30212 35588 30222
rect 35532 30118 35588 30156
rect 34860 30100 34916 30110
rect 34524 29988 34580 29998
rect 34860 29988 34916 30044
rect 34524 29986 34916 29988
rect 34524 29934 34526 29986
rect 34578 29934 34916 29986
rect 34524 29932 34916 29934
rect 34524 29922 34580 29932
rect 35756 29764 35812 31052
rect 35868 31042 35924 31052
rect 36652 30772 36708 30782
rect 35868 30770 36708 30772
rect 35868 30718 36654 30770
rect 36706 30718 36708 30770
rect 35868 30716 36708 30718
rect 35868 30098 35924 30716
rect 36652 30706 36708 30716
rect 36204 30324 36260 30334
rect 36204 30230 36260 30268
rect 36988 30324 37044 33294
rect 37100 33292 37324 33348
rect 37100 31948 37156 33292
rect 37324 33282 37380 33292
rect 37996 33122 38052 36092
rect 38108 34356 38164 34366
rect 38220 34356 38276 39452
rect 38164 34300 38276 34356
rect 38108 34262 38164 34300
rect 37996 33070 37998 33122
rect 38050 33070 38052 33122
rect 37436 32788 37492 32798
rect 37996 32788 38052 33070
rect 37436 32786 38052 32788
rect 37436 32734 37438 32786
rect 37490 32734 38052 32786
rect 37436 32732 38052 32734
rect 38108 33570 38164 33582
rect 38108 33518 38110 33570
rect 38162 33518 38164 33570
rect 38108 32786 38164 33518
rect 38220 33460 38276 33470
rect 38332 33460 38388 39564
rect 38556 39554 38612 39564
rect 38556 37380 38612 37390
rect 38556 37286 38612 37324
rect 38780 36370 38836 36382
rect 38780 36318 38782 36370
rect 38834 36318 38836 36370
rect 38780 35924 38836 36318
rect 38892 36148 38948 41692
rect 39116 41300 39172 41310
rect 39564 41300 39620 42476
rect 39676 42196 39732 42206
rect 39676 41858 39732 42140
rect 40236 42196 40292 42702
rect 39676 41806 39678 41858
rect 39730 41806 39732 41858
rect 39676 41794 39732 41806
rect 39788 41970 39844 41982
rect 39788 41918 39790 41970
rect 39842 41918 39844 41970
rect 39116 41298 39620 41300
rect 39116 41246 39118 41298
rect 39170 41246 39620 41298
rect 39116 41244 39620 41246
rect 39116 41234 39172 41244
rect 39564 40964 39620 40974
rect 39004 40572 39284 40628
rect 39004 40514 39060 40572
rect 39004 40462 39006 40514
rect 39058 40462 39060 40514
rect 39004 40450 39060 40462
rect 39116 40402 39172 40414
rect 39116 40350 39118 40402
rect 39170 40350 39172 40402
rect 39116 39732 39172 40350
rect 39116 39618 39172 39676
rect 39116 39566 39118 39618
rect 39170 39566 39172 39618
rect 39116 39554 39172 39566
rect 39228 40180 39284 40572
rect 39452 40516 39508 40526
rect 39452 40422 39508 40460
rect 39564 40404 39620 40908
rect 39788 40516 39844 41918
rect 39900 41748 39956 41758
rect 39900 41654 39956 41692
rect 39788 40450 39844 40460
rect 39564 40338 39620 40348
rect 39228 39506 39284 40124
rect 39228 39454 39230 39506
rect 39282 39454 39284 39506
rect 39228 39442 39284 39454
rect 39564 39730 39620 39742
rect 39564 39678 39566 39730
rect 39618 39678 39620 39730
rect 39564 39396 39620 39678
rect 40236 39508 40292 42140
rect 40908 41748 40964 44940
rect 41020 44930 41076 44940
rect 41244 44996 41300 45054
rect 41244 44930 41300 44940
rect 41356 44212 41412 46622
rect 41804 46676 41860 46686
rect 41804 45220 41860 46620
rect 41916 45220 41972 45230
rect 41804 45218 41972 45220
rect 41804 45166 41918 45218
rect 41970 45166 41972 45218
rect 41804 45164 41972 45166
rect 41916 45154 41972 45164
rect 41356 44146 41412 44156
rect 41916 44212 41972 44222
rect 41020 44100 41076 44110
rect 41020 43652 41076 44044
rect 41020 43650 41636 43652
rect 41020 43598 41022 43650
rect 41074 43598 41636 43650
rect 41020 43596 41636 43598
rect 41020 43586 41076 43596
rect 41356 42642 41412 42654
rect 41356 42590 41358 42642
rect 41410 42590 41412 42642
rect 41244 42420 41300 42430
rect 41020 41748 41076 41758
rect 40908 41692 41020 41748
rect 41020 41682 41076 41692
rect 41244 40514 41300 42364
rect 41244 40462 41246 40514
rect 41298 40462 41300 40514
rect 40684 40068 40740 40078
rect 39564 39330 39620 39340
rect 39788 39506 40292 39508
rect 39788 39454 40238 39506
rect 40290 39454 40292 39506
rect 39788 39452 40292 39454
rect 39788 39060 39844 39452
rect 40236 39442 40292 39452
rect 40572 39618 40628 39630
rect 40572 39566 40574 39618
rect 40626 39566 40628 39618
rect 40572 39396 40628 39566
rect 40572 39330 40628 39340
rect 39788 38966 39844 39004
rect 39340 37380 39396 37390
rect 39788 37380 39844 37390
rect 39396 37324 39508 37380
rect 39340 37286 39396 37324
rect 39228 37266 39284 37278
rect 39228 37214 39230 37266
rect 39282 37214 39284 37266
rect 39116 36484 39172 36494
rect 39228 36484 39284 37214
rect 39452 36594 39508 37324
rect 39564 37268 39620 37278
rect 39564 37174 39620 37212
rect 39788 37266 39844 37324
rect 39788 37214 39790 37266
rect 39842 37214 39844 37266
rect 39788 37202 39844 37214
rect 40012 37156 40068 37166
rect 40012 37062 40068 37100
rect 39452 36542 39454 36594
rect 39506 36542 39508 36594
rect 39452 36530 39508 36542
rect 39900 37044 39956 37054
rect 39172 36428 39284 36484
rect 39116 36390 39172 36428
rect 39900 36370 39956 36988
rect 40124 37042 40180 37054
rect 40124 36990 40126 37042
rect 40178 36990 40180 37042
rect 39900 36318 39902 36370
rect 39954 36318 39956 36370
rect 39900 36306 39956 36318
rect 40012 36708 40068 36718
rect 38892 36082 38948 36092
rect 38780 35858 38836 35868
rect 39676 35924 39732 35934
rect 39676 35830 39732 35868
rect 40012 35922 40068 36652
rect 40124 36484 40180 36990
rect 40124 36418 40180 36428
rect 40012 35870 40014 35922
rect 40066 35870 40068 35922
rect 40012 35028 40068 35870
rect 40012 34962 40068 34972
rect 40684 35026 40740 40012
rect 41244 40068 41300 40462
rect 41356 40516 41412 42590
rect 41468 42194 41524 43596
rect 41580 43428 41636 43596
rect 41580 43426 41860 43428
rect 41580 43374 41582 43426
rect 41634 43374 41860 43426
rect 41580 43372 41860 43374
rect 41580 43362 41636 43372
rect 41804 42866 41860 43372
rect 41804 42814 41806 42866
rect 41858 42814 41860 42866
rect 41804 42802 41860 42814
rect 41468 42142 41470 42194
rect 41522 42142 41524 42194
rect 41468 42130 41524 42142
rect 41356 40450 41412 40460
rect 41580 40404 41636 40414
rect 41580 40310 41636 40348
rect 41244 40002 41300 40012
rect 40684 34974 40686 35026
rect 40738 34974 40740 35026
rect 40684 34962 40740 34974
rect 40796 39956 40852 39966
rect 40796 35028 40852 39900
rect 41916 39956 41972 44156
rect 42028 43764 42084 46732
rect 42140 46562 42196 47292
rect 42924 46788 42980 46798
rect 43036 46788 43092 48748
rect 42924 46786 43092 46788
rect 42924 46734 42926 46786
rect 42978 46734 43092 46786
rect 42924 46732 43092 46734
rect 43148 48356 43204 48366
rect 42924 46722 42980 46732
rect 42588 46676 42644 46686
rect 42588 46582 42644 46620
rect 43148 46674 43204 48300
rect 43372 47124 43428 49308
rect 44268 49250 44324 50876
rect 44940 50708 44996 52108
rect 45724 52052 45780 52062
rect 45612 52050 45780 52052
rect 45612 51998 45726 52050
rect 45778 51998 45780 52050
rect 45612 51996 45780 51998
rect 45500 51268 45556 51278
rect 45612 51268 45668 51996
rect 45724 51986 45780 51996
rect 45836 51938 45892 51950
rect 45836 51886 45838 51938
rect 45890 51886 45892 51938
rect 45724 51380 45780 51390
rect 45836 51380 45892 51886
rect 46060 51938 46116 51950
rect 46060 51886 46062 51938
rect 46114 51886 46116 51938
rect 46060 51492 46116 51886
rect 46060 51426 46116 51436
rect 46172 51492 46228 51502
rect 46396 51492 46452 53454
rect 47068 52948 47124 53676
rect 47180 53638 47236 53676
rect 47180 52948 47236 52958
rect 47068 52946 47236 52948
rect 47068 52894 47182 52946
rect 47234 52894 47236 52946
rect 47068 52892 47236 52894
rect 47180 52882 47236 52892
rect 47404 52946 47460 53900
rect 47852 53842 47908 53854
rect 48748 53844 48804 55246
rect 49084 55076 49140 55086
rect 49084 54626 49140 55020
rect 49084 54574 49086 54626
rect 49138 54574 49140 54626
rect 49084 54562 49140 54574
rect 49308 54626 49364 54638
rect 49308 54574 49310 54626
rect 49362 54574 49364 54626
rect 49308 54516 49364 54574
rect 49308 54450 49364 54460
rect 47852 53790 47854 53842
rect 47906 53790 47908 53842
rect 47852 53732 47908 53790
rect 48636 53788 48804 53844
rect 49196 54402 49252 54414
rect 49196 54350 49198 54402
rect 49250 54350 49252 54402
rect 47852 53666 47908 53676
rect 47964 53730 48020 53742
rect 47964 53678 47966 53730
rect 48018 53678 48020 53730
rect 47404 52894 47406 52946
rect 47458 52894 47460 52946
rect 47404 52882 47460 52894
rect 47628 52724 47684 52734
rect 47516 52722 47908 52724
rect 47516 52670 47630 52722
rect 47682 52670 47908 52722
rect 47516 52668 47908 52670
rect 47516 51940 47572 52668
rect 47628 52658 47684 52668
rect 47292 51884 47572 51940
rect 47628 52050 47684 52062
rect 47628 51998 47630 52050
rect 47682 51998 47684 52050
rect 47292 51602 47348 51884
rect 47292 51550 47294 51602
rect 47346 51550 47348 51602
rect 47292 51538 47348 51550
rect 46172 51490 46452 51492
rect 46172 51438 46174 51490
rect 46226 51438 46452 51490
rect 46172 51436 46452 51438
rect 46844 51492 46900 51502
rect 46172 51426 46228 51436
rect 45724 51378 45892 51380
rect 45724 51326 45726 51378
rect 45778 51326 45892 51378
rect 45724 51324 45892 51326
rect 45724 51314 45780 51324
rect 45500 51266 45668 51268
rect 45500 51214 45502 51266
rect 45554 51214 45668 51266
rect 45500 51212 45668 51214
rect 45500 50932 45556 51212
rect 45500 50866 45556 50876
rect 44940 50706 45108 50708
rect 44940 50654 44942 50706
rect 44994 50654 45108 50706
rect 44940 50652 45108 50654
rect 44940 50642 44996 50652
rect 44380 50482 44436 50494
rect 44380 50430 44382 50482
rect 44434 50430 44436 50482
rect 44380 50428 44436 50430
rect 44380 50372 44548 50428
rect 44492 50306 44548 50316
rect 45052 49922 45108 50652
rect 45164 50594 45220 50606
rect 45164 50542 45166 50594
rect 45218 50542 45220 50594
rect 45164 50484 45220 50542
rect 45220 50428 45444 50484
rect 45164 50418 45220 50428
rect 45052 49870 45054 49922
rect 45106 49870 45108 49922
rect 45052 49858 45108 49870
rect 45388 49810 45444 50428
rect 45836 50482 45892 51324
rect 45836 50430 45838 50482
rect 45890 50430 45892 50482
rect 45836 50428 45892 50430
rect 46620 50594 46676 50606
rect 46620 50542 46622 50594
rect 46674 50542 46676 50594
rect 46620 50484 46676 50542
rect 46844 50594 46900 51436
rect 47404 51492 47460 51502
rect 47404 51398 47460 51436
rect 46844 50542 46846 50594
rect 46898 50542 46900 50594
rect 46844 50530 46900 50542
rect 46956 51378 47012 51390
rect 46956 51326 46958 51378
rect 47010 51326 47012 51378
rect 46956 50482 47012 51326
rect 46956 50430 46958 50482
rect 47010 50430 47012 50482
rect 46956 50428 47012 50430
rect 45836 50372 46004 50428
rect 45388 49758 45390 49810
rect 45442 49758 45444 49810
rect 45388 49746 45444 49758
rect 45948 49810 46004 50372
rect 45948 49758 45950 49810
rect 46002 49758 46004 49810
rect 45948 49746 46004 49758
rect 46508 50372 46676 50428
rect 46844 50372 47012 50428
rect 47068 51378 47124 51390
rect 47068 51326 47070 51378
rect 47122 51326 47124 51378
rect 47068 50484 47124 51326
rect 47628 50932 47684 51998
rect 47852 52050 47908 52668
rect 47964 52386 48020 53678
rect 48636 53396 48692 53788
rect 48748 53620 48804 53630
rect 49084 53620 49140 53630
rect 48748 53618 49140 53620
rect 48748 53566 48750 53618
rect 48802 53566 49086 53618
rect 49138 53566 49140 53618
rect 48748 53564 49140 53566
rect 48748 53554 48804 53564
rect 49084 53554 49140 53564
rect 48636 53340 48804 53396
rect 47964 52334 47966 52386
rect 48018 52334 48020 52386
rect 47964 52322 48020 52334
rect 48076 52722 48132 52734
rect 48076 52670 48078 52722
rect 48130 52670 48132 52722
rect 47852 51998 47854 52050
rect 47906 51998 47908 52050
rect 47852 51986 47908 51998
rect 47404 50876 47908 50932
rect 47404 50818 47460 50876
rect 47404 50766 47406 50818
rect 47458 50766 47460 50818
rect 47404 50754 47460 50766
rect 47740 50596 47796 50606
rect 47068 50418 47124 50428
rect 47516 50594 47796 50596
rect 47516 50542 47742 50594
rect 47794 50542 47796 50594
rect 47516 50540 47796 50542
rect 46060 49698 46116 49710
rect 46060 49646 46062 49698
rect 46114 49646 46116 49698
rect 45388 49588 45444 49598
rect 45388 49494 45444 49532
rect 44268 49198 44270 49250
rect 44322 49198 44324 49250
rect 44268 49186 44324 49198
rect 43596 49140 43652 49150
rect 43596 49046 43652 49084
rect 45948 49028 46004 49038
rect 46060 49028 46116 49646
rect 45724 49026 46116 49028
rect 45724 48974 45950 49026
rect 46002 48974 46116 49026
rect 45724 48972 46116 48974
rect 46172 49588 46228 49598
rect 46172 49026 46228 49532
rect 46172 48974 46174 49026
rect 46226 48974 46228 49026
rect 43932 48916 43988 48926
rect 43932 48822 43988 48860
rect 43484 48804 43540 48814
rect 43596 48804 43652 48814
rect 43484 48802 43596 48804
rect 43484 48750 43486 48802
rect 43538 48750 43596 48802
rect 43484 48748 43596 48750
rect 43484 48738 43540 48748
rect 43484 47124 43540 47134
rect 43372 47068 43484 47124
rect 43484 47058 43540 47068
rect 43148 46622 43150 46674
rect 43202 46622 43204 46674
rect 43148 46610 43204 46622
rect 42140 46510 42142 46562
rect 42194 46510 42196 46562
rect 42140 46498 42196 46510
rect 42700 45332 42756 45342
rect 42252 45108 42308 45118
rect 42252 45014 42308 45052
rect 42476 45106 42532 45118
rect 42476 45054 42478 45106
rect 42530 45054 42532 45106
rect 42364 44996 42420 45006
rect 42364 44902 42420 44940
rect 42364 44322 42420 44334
rect 42364 44270 42366 44322
rect 42418 44270 42420 44322
rect 42028 43708 42196 43764
rect 42028 43538 42084 43550
rect 42028 43486 42030 43538
rect 42082 43486 42084 43538
rect 42028 42756 42084 43486
rect 42028 42662 42084 42700
rect 42140 42420 42196 43708
rect 42364 43652 42420 44270
rect 42476 44212 42532 45054
rect 42700 44434 42756 45276
rect 42700 44382 42702 44434
rect 42754 44382 42756 44434
rect 42700 44370 42756 44382
rect 43484 44324 43540 44334
rect 43596 44324 43652 48748
rect 44156 48804 44212 48814
rect 44156 48710 44212 48748
rect 43932 48580 43988 48590
rect 43932 48242 43988 48524
rect 44940 48468 44996 48478
rect 44940 48374 44996 48412
rect 44044 48356 44100 48366
rect 44044 48262 44100 48300
rect 44604 48356 44660 48366
rect 43932 48190 43934 48242
rect 43986 48190 43988 48242
rect 43932 48178 43988 48190
rect 44156 46788 44212 46798
rect 44156 46694 44212 46732
rect 43932 46674 43988 46686
rect 43932 46622 43934 46674
rect 43986 46622 43988 46674
rect 43820 45892 43876 45902
rect 43820 45798 43876 45836
rect 43708 45780 43764 45790
rect 43708 45686 43764 45724
rect 43484 44322 43652 44324
rect 43484 44270 43486 44322
rect 43538 44270 43652 44322
rect 43484 44268 43652 44270
rect 43484 44258 43540 44268
rect 42700 44212 42756 44222
rect 42476 44156 42700 44212
rect 42756 44156 43092 44212
rect 42700 44118 42756 44156
rect 43036 43762 43092 44156
rect 43036 43710 43038 43762
rect 43090 43710 43092 43762
rect 43036 43698 43092 43710
rect 42812 43652 42868 43662
rect 42364 43650 42868 43652
rect 42364 43598 42814 43650
rect 42866 43598 42868 43650
rect 42364 43596 42868 43598
rect 42364 43426 42420 43596
rect 42812 43586 42868 43596
rect 42364 43374 42366 43426
rect 42418 43374 42420 43426
rect 42364 43362 42420 43374
rect 43148 43316 43204 43326
rect 43148 43222 43204 43260
rect 43148 42868 43204 42878
rect 43148 42774 43204 42812
rect 42700 42644 42756 42654
rect 43036 42644 43092 42654
rect 42700 42642 43092 42644
rect 42700 42590 42702 42642
rect 42754 42590 43038 42642
rect 43090 42590 43092 42642
rect 42700 42588 43092 42590
rect 42700 42578 42756 42588
rect 43036 42578 43092 42588
rect 42140 42354 42196 42364
rect 43260 42530 43316 42542
rect 43260 42478 43262 42530
rect 43314 42478 43316 42530
rect 43260 42420 43316 42478
rect 43260 42354 43316 42364
rect 43484 42530 43540 42542
rect 43484 42478 43486 42530
rect 43538 42478 43540 42530
rect 42476 41748 42532 41758
rect 41916 39890 41972 39900
rect 42028 40516 42084 40526
rect 41132 39620 41188 39630
rect 41580 39620 41636 39630
rect 41132 39618 41636 39620
rect 41132 39566 41134 39618
rect 41186 39566 41582 39618
rect 41634 39566 41636 39618
rect 41132 39564 41636 39566
rect 41132 39554 41188 39564
rect 41580 39554 41636 39564
rect 41804 39620 41860 39630
rect 41020 39394 41076 39406
rect 41020 39342 41022 39394
rect 41074 39342 41076 39394
rect 41020 38668 41076 39342
rect 41468 39396 41524 39406
rect 41692 39396 41748 39406
rect 41468 39302 41524 39340
rect 41580 39394 41748 39396
rect 41580 39342 41694 39394
rect 41746 39342 41748 39394
rect 41580 39340 41748 39342
rect 41244 39060 41300 39070
rect 41580 39060 41636 39340
rect 41692 39330 41748 39340
rect 41300 39004 41636 39060
rect 41692 39060 41748 39070
rect 41804 39060 41860 39564
rect 41692 39058 41860 39060
rect 41692 39006 41694 39058
rect 41746 39006 41860 39058
rect 41692 39004 41860 39006
rect 42028 39060 42084 40460
rect 42476 40402 42532 41692
rect 42476 40350 42478 40402
rect 42530 40350 42532 40402
rect 42476 40338 42532 40350
rect 43484 40626 43540 42478
rect 43484 40574 43486 40626
rect 43538 40574 43540 40626
rect 43148 40292 43204 40302
rect 43148 40290 43428 40292
rect 43148 40238 43150 40290
rect 43202 40238 43428 40290
rect 43148 40236 43428 40238
rect 43148 40226 43204 40236
rect 43148 40068 43204 40078
rect 43148 39732 43204 40012
rect 42700 39676 43204 39732
rect 42140 39620 42196 39630
rect 42364 39620 42420 39630
rect 42196 39618 42420 39620
rect 42196 39566 42366 39618
rect 42418 39566 42420 39618
rect 42196 39564 42420 39566
rect 42140 39526 42196 39564
rect 42364 39554 42420 39564
rect 42700 39508 42756 39676
rect 43148 39618 43204 39676
rect 43148 39566 43150 39618
rect 43202 39566 43204 39618
rect 43148 39554 43204 39566
rect 43372 39618 43428 40236
rect 43484 40068 43540 40574
rect 43484 40002 43540 40012
rect 43372 39566 43374 39618
rect 43426 39566 43428 39618
rect 42476 39506 42756 39508
rect 42476 39454 42702 39506
rect 42754 39454 42756 39506
rect 42476 39452 42756 39454
rect 42140 39060 42196 39070
rect 42028 39058 42196 39060
rect 42028 39006 42142 39058
rect 42194 39006 42196 39058
rect 42028 39004 42196 39006
rect 41244 38966 41300 39004
rect 41692 38994 41748 39004
rect 42140 38994 42196 39004
rect 42252 38948 42308 38958
rect 42476 38948 42532 39452
rect 42700 39442 42756 39452
rect 42252 38946 42532 38948
rect 42252 38894 42254 38946
rect 42306 38894 42532 38946
rect 42252 38892 42532 38894
rect 42812 39396 42868 39406
rect 42252 38882 42308 38892
rect 41580 38836 41636 38846
rect 41580 38722 41636 38780
rect 41580 38670 41582 38722
rect 41634 38670 41636 38722
rect 41020 38612 41188 38668
rect 41580 38658 41636 38670
rect 41132 37378 41188 38612
rect 42140 38612 42196 38622
rect 42140 38518 42196 38556
rect 42812 38050 42868 39340
rect 43372 39284 43428 39566
rect 43148 39228 43428 39284
rect 43484 39844 43540 39854
rect 43484 39618 43540 39788
rect 43484 39566 43486 39618
rect 43538 39566 43540 39618
rect 43036 38948 43092 38958
rect 42812 37998 42814 38050
rect 42866 37998 42868 38050
rect 42812 37986 42868 37998
rect 42924 38892 43036 38948
rect 42476 37940 42532 37950
rect 42476 37846 42532 37884
rect 42588 37826 42644 37838
rect 42588 37774 42590 37826
rect 42642 37774 42644 37826
rect 41916 37492 41972 37502
rect 41916 37398 41972 37436
rect 41132 37326 41134 37378
rect 41186 37326 41188 37378
rect 40908 37268 40964 37278
rect 40908 37174 40964 37212
rect 41132 37044 41188 37326
rect 41804 37266 41860 37278
rect 41804 37214 41806 37266
rect 41858 37214 41860 37266
rect 41804 37156 41860 37214
rect 41804 37090 41860 37100
rect 41132 36978 41188 36988
rect 42588 36708 42644 37774
rect 42812 36932 42868 36942
rect 42028 36652 42756 36708
rect 40908 36484 40964 36494
rect 40908 36390 40964 36428
rect 41580 36372 41636 36382
rect 41580 36278 41636 36316
rect 41916 36370 41972 36382
rect 41916 36318 41918 36370
rect 41970 36318 41972 36370
rect 41916 36036 41972 36318
rect 41916 35970 41972 35980
rect 42028 36370 42084 36652
rect 42252 36484 42308 36494
rect 42588 36484 42644 36494
rect 42252 36482 42644 36484
rect 42252 36430 42254 36482
rect 42306 36430 42590 36482
rect 42642 36430 42644 36482
rect 42252 36428 42644 36430
rect 42252 36418 42308 36428
rect 42588 36418 42644 36428
rect 42028 36318 42030 36370
rect 42082 36318 42084 36370
rect 42028 35924 42084 36318
rect 42028 35858 42084 35868
rect 42700 35922 42756 36652
rect 42812 36484 42868 36876
rect 42812 36390 42868 36428
rect 42700 35870 42702 35922
rect 42754 35870 42756 35922
rect 42700 35858 42756 35870
rect 40796 34972 41524 35028
rect 40348 34914 40404 34926
rect 40348 34862 40350 34914
rect 40402 34862 40404 34914
rect 40012 34804 40068 34814
rect 39116 34132 39172 34142
rect 39116 34038 39172 34076
rect 39788 34132 39844 34142
rect 39788 34038 39844 34076
rect 38276 33404 38388 33460
rect 38668 34020 38724 34030
rect 38220 33394 38276 33404
rect 38668 33236 38724 33964
rect 38108 32734 38110 32786
rect 38162 32734 38164 32786
rect 37436 32722 37492 32732
rect 38108 32722 38164 32734
rect 38556 33180 38724 33236
rect 39452 34018 39508 34030
rect 39452 33966 39454 34018
rect 39506 33966 39508 34018
rect 37212 32676 37268 32686
rect 37212 32582 37268 32620
rect 38332 32676 38388 32686
rect 38332 32582 38388 32620
rect 37884 32562 37940 32574
rect 37884 32510 37886 32562
rect 37938 32510 37940 32562
rect 37324 32452 37380 32462
rect 37884 32452 37940 32510
rect 38220 32564 38276 32574
rect 38220 32470 38276 32508
rect 37324 32450 37716 32452
rect 37324 32398 37326 32450
rect 37378 32398 37716 32450
rect 37324 32396 37716 32398
rect 37324 32386 37380 32396
rect 37660 31948 37716 32396
rect 37884 32386 37940 32396
rect 38556 32116 38612 33180
rect 38780 33124 38836 33134
rect 38668 33122 38836 33124
rect 38668 33070 38782 33122
rect 38834 33070 38836 33122
rect 38668 33068 38836 33070
rect 38668 32788 38724 33068
rect 38780 33058 38836 33068
rect 39452 33012 39508 33966
rect 40012 33346 40068 34748
rect 40348 34132 40404 34862
rect 41356 34802 41412 34814
rect 41356 34750 41358 34802
rect 41410 34750 41412 34802
rect 41020 34692 41076 34702
rect 40348 34066 40404 34076
rect 40908 34690 41076 34692
rect 40908 34638 41022 34690
rect 41074 34638 41076 34690
rect 40908 34636 41076 34638
rect 40908 34130 40964 34636
rect 41020 34626 41076 34636
rect 40908 34078 40910 34130
rect 40962 34078 40964 34130
rect 40908 34020 40964 34078
rect 41132 34132 41188 34142
rect 41132 34038 41188 34076
rect 40908 33954 40964 33964
rect 40012 33294 40014 33346
rect 40066 33294 40068 33346
rect 40012 33282 40068 33294
rect 40348 33236 40404 33246
rect 40348 33142 40404 33180
rect 41356 33236 41412 34750
rect 41468 34354 41524 34972
rect 41468 34302 41470 34354
rect 41522 34302 41524 34354
rect 41468 34290 41524 34302
rect 41356 33170 41412 33180
rect 42140 33346 42196 33358
rect 42924 33348 42980 38892
rect 43036 38854 43092 38892
rect 43148 38834 43204 39228
rect 43148 38782 43150 38834
rect 43202 38782 43204 38834
rect 43148 38770 43204 38782
rect 43484 38834 43540 39566
rect 43484 38782 43486 38834
rect 43538 38782 43540 38834
rect 43484 38770 43540 38782
rect 43596 38836 43652 44268
rect 43820 42532 43876 42542
rect 43820 41970 43876 42476
rect 43932 42084 43988 46622
rect 44604 46564 44660 48300
rect 45612 48354 45668 48366
rect 45612 48302 45614 48354
rect 45666 48302 45668 48354
rect 44940 48244 44996 48254
rect 44268 46562 44660 46564
rect 44268 46510 44606 46562
rect 44658 46510 44660 46562
rect 44268 46508 44660 46510
rect 44268 46452 44324 46508
rect 44604 46498 44660 46508
rect 44828 48188 44940 48244
rect 44044 46396 44324 46452
rect 44044 45890 44100 46396
rect 44044 45838 44046 45890
rect 44098 45838 44100 45890
rect 44044 45826 44100 45838
rect 44268 45778 44324 45790
rect 44268 45726 44270 45778
rect 44322 45726 44324 45778
rect 44156 45556 44212 45566
rect 43932 42028 44100 42084
rect 43820 41918 43822 41970
rect 43874 41918 43876 41970
rect 43820 41906 43876 41918
rect 43932 41858 43988 41870
rect 43932 41806 43934 41858
rect 43986 41806 43988 41858
rect 43932 40628 43988 41806
rect 43820 40572 43988 40628
rect 43820 40292 43876 40572
rect 43820 39396 43876 40236
rect 44044 40402 44100 42028
rect 44044 40350 44046 40402
rect 44098 40350 44100 40402
rect 43932 39620 43988 39630
rect 43932 39526 43988 39564
rect 43820 39330 43876 39340
rect 44044 38948 44100 40350
rect 44044 38882 44100 38892
rect 43596 38770 43652 38780
rect 43260 38724 43316 38762
rect 43260 38658 43316 38668
rect 43932 38612 43988 38622
rect 43932 37490 43988 38556
rect 43932 37438 43934 37490
rect 43986 37438 43988 37490
rect 43708 37266 43764 37278
rect 43708 37214 43710 37266
rect 43762 37214 43764 37266
rect 43484 36372 43540 36382
rect 43708 36372 43764 37214
rect 43820 37154 43876 37166
rect 43820 37102 43822 37154
rect 43874 37102 43876 37154
rect 43820 36596 43876 37102
rect 43820 36530 43876 36540
rect 43484 36370 43764 36372
rect 43484 36318 43486 36370
rect 43538 36318 43764 36370
rect 43484 36316 43764 36318
rect 43820 36370 43876 36382
rect 43820 36318 43822 36370
rect 43874 36318 43876 36370
rect 43036 36260 43092 36270
rect 43036 35924 43092 36204
rect 43036 35922 43428 35924
rect 43036 35870 43038 35922
rect 43090 35870 43428 35922
rect 43036 35868 43428 35870
rect 43036 35858 43092 35868
rect 43372 34354 43428 35868
rect 43484 35700 43540 36316
rect 43708 36036 43764 36046
rect 43820 36036 43876 36318
rect 43764 35980 43876 36036
rect 43708 35970 43764 35980
rect 43596 35700 43652 35710
rect 43484 35698 43652 35700
rect 43484 35646 43598 35698
rect 43650 35646 43652 35698
rect 43484 35644 43652 35646
rect 43596 35634 43652 35644
rect 43932 35698 43988 37438
rect 44044 36484 44100 36494
rect 44044 36390 44100 36428
rect 44156 36260 44212 45500
rect 44268 45108 44324 45726
rect 44828 45332 44884 48188
rect 44940 48150 44996 48188
rect 45612 48244 45668 48302
rect 45612 48178 45668 48188
rect 45724 48130 45780 48972
rect 45948 48962 46004 48972
rect 46172 48962 46228 48974
rect 46508 49026 46564 50372
rect 46844 49922 46900 50372
rect 47516 50034 47572 50540
rect 47740 50530 47796 50540
rect 47516 49982 47518 50034
rect 47570 49982 47572 50034
rect 47516 49970 47572 49982
rect 46844 49870 46846 49922
rect 46898 49870 46900 49922
rect 46844 49858 46900 49870
rect 47852 49922 47908 50876
rect 47852 49870 47854 49922
rect 47906 49870 47908 49922
rect 47852 49858 47908 49870
rect 47964 50596 48020 50606
rect 46508 48974 46510 49026
rect 46562 48974 46564 49026
rect 46508 48962 46564 48974
rect 47180 49810 47236 49822
rect 47180 49758 47182 49810
rect 47234 49758 47236 49810
rect 46060 48804 46116 48814
rect 46060 48710 46116 48748
rect 47180 48804 47236 49758
rect 47628 49810 47684 49822
rect 47628 49758 47630 49810
rect 47682 49758 47684 49810
rect 47628 49140 47684 49758
rect 47852 49252 47908 49262
rect 47964 49252 48020 50540
rect 48076 50482 48132 52670
rect 48636 50596 48692 50606
rect 48636 50502 48692 50540
rect 48076 50430 48078 50482
rect 48130 50430 48132 50482
rect 48076 50418 48132 50430
rect 48748 50428 48804 53340
rect 49196 53060 49252 54350
rect 49532 54068 49588 56028
rect 49644 55412 49700 55422
rect 49644 55318 49700 55356
rect 49980 55076 50036 55086
rect 49980 54514 50036 55020
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 51100 54852 51156 59200
rect 52220 56308 52276 56318
rect 52220 56214 52276 56252
rect 51212 56084 51268 56094
rect 51212 55990 51268 56028
rect 52444 55412 52500 59200
rect 53116 56308 53172 59200
rect 53788 56642 53844 59200
rect 53788 56590 53790 56642
rect 53842 56590 53844 56642
rect 53788 56578 53844 56590
rect 53116 56242 53172 56252
rect 54124 56308 54180 56318
rect 54124 56214 54180 56252
rect 54460 56308 54516 59200
rect 54460 56242 54516 56252
rect 55020 56642 55076 56654
rect 55020 56590 55022 56642
rect 55074 56590 55076 56642
rect 55020 56306 55076 56590
rect 55020 56254 55022 56306
rect 55074 56254 55076 56306
rect 55020 56242 55076 56254
rect 55132 55972 55188 59200
rect 55468 56308 55524 56318
rect 55468 56214 55524 56252
rect 55132 55906 55188 55916
rect 55916 55972 55972 55982
rect 55916 55878 55972 55916
rect 58156 55860 58212 55870
rect 58156 55766 58212 55804
rect 52444 55346 52500 55356
rect 53676 55412 53732 55422
rect 53676 55318 53732 55356
rect 51772 55300 51828 55310
rect 51100 54786 51156 54796
rect 51436 55298 51828 55300
rect 51436 55246 51774 55298
rect 51826 55246 51828 55298
rect 51436 55244 51828 55246
rect 50876 54628 50932 54638
rect 51436 54628 51492 55244
rect 51772 55234 51828 55244
rect 53004 55298 53060 55310
rect 53004 55246 53006 55298
rect 53058 55246 53060 55298
rect 50876 54626 51492 54628
rect 50876 54574 50878 54626
rect 50930 54574 51492 54626
rect 50876 54572 51492 54574
rect 51548 55074 51604 55086
rect 51548 55022 51550 55074
rect 51602 55022 51604 55074
rect 50876 54562 50932 54572
rect 49980 54462 49982 54514
rect 50034 54462 50036 54514
rect 49980 54450 50036 54462
rect 50092 54516 50148 54526
rect 49420 54012 49588 54068
rect 49420 53618 49476 54012
rect 49420 53566 49422 53618
rect 49474 53566 49476 53618
rect 49420 53554 49476 53566
rect 49644 53730 49700 53742
rect 49644 53678 49646 53730
rect 49698 53678 49700 53730
rect 49644 53620 49700 53678
rect 50092 53732 50148 54460
rect 51548 54514 51604 55022
rect 52332 54852 52388 54862
rect 52332 54738 52388 54796
rect 52332 54686 52334 54738
rect 52386 54686 52388 54738
rect 52332 54674 52388 54686
rect 51548 54462 51550 54514
rect 51602 54462 51604 54514
rect 51548 54450 51604 54462
rect 50204 54402 50260 54414
rect 50204 54350 50206 54402
rect 50258 54350 50260 54402
rect 50204 53842 50260 54350
rect 50204 53790 50206 53842
rect 50258 53790 50260 53842
rect 50204 53778 50260 53790
rect 50876 54180 50932 54190
rect 50092 53638 50148 53676
rect 49644 53554 49700 53564
rect 50316 53508 50372 53518
rect 50316 53414 50372 53452
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 49196 52994 49252 53004
rect 50652 53060 50708 53070
rect 50652 52966 50708 53004
rect 50876 52834 50932 54124
rect 51324 53842 51380 53854
rect 51324 53790 51326 53842
rect 51378 53790 51380 53842
rect 50988 53732 51044 53742
rect 50988 53638 51044 53676
rect 51324 53508 51380 53790
rect 51660 53620 51716 53630
rect 51660 53526 51716 53564
rect 52668 53620 52724 53630
rect 52668 53526 52724 53564
rect 53004 53618 53060 55246
rect 57708 55188 57764 55198
rect 57708 55094 57764 55132
rect 58156 55074 58212 55086
rect 58156 55022 58158 55074
rect 58210 55022 58212 55074
rect 58156 54516 58212 55022
rect 58156 54450 58212 54460
rect 53004 53566 53006 53618
rect 53058 53566 53060 53618
rect 53004 53554 53060 53566
rect 50876 52782 50878 52834
rect 50930 52782 50932 52834
rect 50876 52770 50932 52782
rect 50988 52946 51044 52958
rect 50988 52894 50990 52946
rect 51042 52894 51044 52946
rect 50988 51938 51044 52894
rect 51324 52274 51380 53452
rect 58156 53058 58212 53070
rect 58156 53006 58158 53058
rect 58210 53006 58212 53058
rect 51772 52946 51828 52958
rect 51772 52894 51774 52946
rect 51826 52894 51828 52946
rect 51324 52222 51326 52274
rect 51378 52222 51380 52274
rect 51324 52210 51380 52222
rect 51660 52834 51716 52846
rect 51660 52782 51662 52834
rect 51714 52782 51716 52834
rect 51436 52164 51492 52202
rect 51660 52164 51716 52782
rect 51492 52108 51716 52164
rect 51772 52274 51828 52894
rect 58156 52500 58212 53006
rect 58156 52434 58212 52444
rect 51772 52222 51774 52274
rect 51826 52222 51828 52274
rect 51436 52098 51492 52108
rect 50988 51886 50990 51938
rect 51042 51886 51044 51938
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50876 51378 50932 51390
rect 50876 51326 50878 51378
rect 50930 51326 50932 51378
rect 50428 51268 50484 51278
rect 50428 50594 50484 51212
rect 50428 50542 50430 50594
rect 50482 50542 50484 50594
rect 50428 50530 50484 50542
rect 50652 50484 50708 50494
rect 48636 50372 48804 50428
rect 50540 50428 50652 50484
rect 50540 50372 50596 50428
rect 50652 50418 50708 50428
rect 50764 50484 50820 50494
rect 50876 50484 50932 51326
rect 50988 50596 51044 51886
rect 51100 52052 51156 52062
rect 51100 51716 51156 51996
rect 51212 51940 51268 51950
rect 51212 51938 51604 51940
rect 51212 51886 51214 51938
rect 51266 51886 51604 51938
rect 51212 51884 51604 51886
rect 51212 51874 51268 51884
rect 51100 51660 51268 51716
rect 50988 50530 51044 50540
rect 51100 51490 51156 51502
rect 51100 51438 51102 51490
rect 51154 51438 51156 51490
rect 50764 50482 50932 50484
rect 50764 50430 50766 50482
rect 50818 50430 50932 50482
rect 50764 50428 50932 50430
rect 50764 50418 50820 50428
rect 48636 50370 48692 50372
rect 48636 50318 48638 50370
rect 48690 50318 48692 50370
rect 48636 50306 48692 50318
rect 50428 50316 50596 50372
rect 50428 50034 50484 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50428 49982 50430 50034
rect 50482 49982 50484 50034
rect 50428 49970 50484 49982
rect 49868 49812 49924 49822
rect 49756 49252 49812 49262
rect 47852 49250 48020 49252
rect 47852 49198 47854 49250
rect 47906 49198 48020 49250
rect 47852 49196 48020 49198
rect 48972 49250 49812 49252
rect 48972 49198 49758 49250
rect 49810 49198 49812 49250
rect 48972 49196 49812 49198
rect 47852 49186 47908 49196
rect 47740 49140 47796 49150
rect 47628 49084 47740 49140
rect 47180 48738 47236 48748
rect 47516 48914 47572 48926
rect 47516 48862 47518 48914
rect 47570 48862 47572 48914
rect 47516 48804 47572 48862
rect 47740 48914 47796 49084
rect 48972 49138 49028 49196
rect 48972 49086 48974 49138
rect 49026 49086 49028 49138
rect 48972 49074 49028 49086
rect 47740 48862 47742 48914
rect 47794 48862 47796 48914
rect 47740 48850 47796 48862
rect 49084 48916 49140 48926
rect 49084 48822 49140 48860
rect 47516 48738 47572 48748
rect 49756 48242 49812 49196
rect 49868 49026 49924 49756
rect 50092 49700 50148 49710
rect 50092 49138 50148 49644
rect 50876 49252 50932 50428
rect 51100 50484 51156 51438
rect 51100 50390 51156 50428
rect 51212 51380 51268 51660
rect 51548 51604 51604 51884
rect 51660 51604 51716 51614
rect 51772 51604 51828 52222
rect 51548 51602 51828 51604
rect 51548 51550 51662 51602
rect 51714 51550 51828 51602
rect 51548 51548 51828 51550
rect 51884 51938 51940 51950
rect 51884 51886 51886 51938
rect 51938 51886 51940 51938
rect 51660 51538 51716 51548
rect 50988 49252 51044 49262
rect 50876 49250 51044 49252
rect 50876 49198 50990 49250
rect 51042 49198 51044 49250
rect 50876 49196 51044 49198
rect 50988 49186 51044 49196
rect 50092 49086 50094 49138
rect 50146 49086 50148 49138
rect 50092 49074 50148 49086
rect 49868 48974 49870 49026
rect 49922 48974 49924 49026
rect 49868 48962 49924 48974
rect 50876 48916 50932 48926
rect 50876 48822 50932 48860
rect 50988 48802 51044 48814
rect 50988 48750 50990 48802
rect 51042 48750 51044 48802
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 49756 48190 49758 48242
rect 49810 48190 49812 48242
rect 49756 48178 49812 48190
rect 49980 48468 50036 48478
rect 49980 48242 50036 48412
rect 50988 48468 51044 48750
rect 50988 48402 51044 48412
rect 49980 48190 49982 48242
rect 50034 48190 50036 48242
rect 49980 48178 50036 48190
rect 45724 48078 45726 48130
rect 45778 48078 45780 48130
rect 45724 48066 45780 48078
rect 50652 48130 50708 48142
rect 50652 48078 50654 48130
rect 50706 48078 50708 48130
rect 45388 48020 45444 48030
rect 45388 47926 45444 47964
rect 46060 47628 46676 47684
rect 45500 47348 45556 47358
rect 45500 47254 45556 47292
rect 45612 47234 45668 47246
rect 45612 47182 45614 47234
rect 45666 47182 45668 47234
rect 45164 47124 45220 47134
rect 45164 46786 45220 47068
rect 45164 46734 45166 46786
rect 45218 46734 45220 46786
rect 45052 46674 45108 46686
rect 45052 46622 45054 46674
rect 45106 46622 45108 46674
rect 45052 46116 45108 46622
rect 45052 46050 45108 46060
rect 44940 45556 44996 45566
rect 45164 45556 45220 46734
rect 45388 46676 45444 46686
rect 45388 45890 45444 46620
rect 45388 45838 45390 45890
rect 45442 45838 45444 45890
rect 45388 45826 45444 45838
rect 45612 46452 45668 47182
rect 46060 46562 46116 47628
rect 46060 46510 46062 46562
rect 46114 46510 46116 46562
rect 46060 46452 46116 46510
rect 45612 46396 46116 46452
rect 46396 47460 46452 47470
rect 46396 46452 46452 47404
rect 46620 47458 46676 47628
rect 49308 47572 49364 47582
rect 49308 47478 49364 47516
rect 50428 47570 50484 47582
rect 50428 47518 50430 47570
rect 50482 47518 50484 47570
rect 46620 47406 46622 47458
rect 46674 47406 46676 47458
rect 46620 47394 46676 47406
rect 49532 47460 49588 47470
rect 49532 47366 49588 47404
rect 50428 47460 50484 47518
rect 50428 47394 50484 47404
rect 50652 47572 50708 48078
rect 50652 47458 50708 47516
rect 50652 47406 50654 47458
rect 50706 47406 50708 47458
rect 50652 47394 50708 47406
rect 46956 47346 47012 47358
rect 46956 47294 46958 47346
rect 47010 47294 47012 47346
rect 46844 47234 46900 47246
rect 46844 47182 46846 47234
rect 46898 47182 46900 47234
rect 46508 46788 46564 46798
rect 46508 46694 46564 46732
rect 46732 46788 46788 46798
rect 46396 46396 46676 46452
rect 45500 45780 45556 45790
rect 45612 45780 45668 46396
rect 45724 45892 45780 45902
rect 46508 45892 46564 45902
rect 45724 45890 46564 45892
rect 45724 45838 45726 45890
rect 45778 45838 46510 45890
rect 46562 45838 46564 45890
rect 45724 45836 46564 45838
rect 45724 45826 45780 45836
rect 46508 45826 46564 45836
rect 45500 45778 45668 45780
rect 45500 45726 45502 45778
rect 45554 45726 45668 45778
rect 45500 45724 45668 45726
rect 45500 45714 45556 45724
rect 46620 45668 46676 46396
rect 46732 45892 46788 46732
rect 46844 46452 46900 47182
rect 46956 46676 47012 47294
rect 49868 47234 49924 47246
rect 49868 47182 49870 47234
rect 49922 47182 49924 47234
rect 47516 46676 47572 46686
rect 47012 46674 47572 46676
rect 47012 46622 47518 46674
rect 47570 46622 47572 46674
rect 47012 46620 47572 46622
rect 46956 46582 47012 46620
rect 47516 46610 47572 46620
rect 49868 46676 49924 47182
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 51100 46788 51156 46798
rect 51212 46788 51268 51324
rect 51548 51378 51604 51390
rect 51548 51326 51550 51378
rect 51602 51326 51604 51378
rect 51548 51268 51604 51326
rect 51548 51202 51604 51212
rect 51660 50596 51716 50606
rect 51660 50502 51716 50540
rect 51884 50484 51940 51886
rect 53900 51490 53956 51502
rect 53900 51438 53902 51490
rect 53954 51438 53956 51490
rect 52332 51380 52388 51390
rect 52332 51266 52388 51324
rect 52332 51214 52334 51266
rect 52386 51214 52388 51266
rect 52332 51202 52388 51214
rect 52780 51378 52836 51390
rect 52780 51326 52782 51378
rect 52834 51326 52836 51378
rect 52780 50818 52836 51326
rect 53228 51380 53284 51390
rect 53564 51380 53620 51390
rect 53228 51378 53620 51380
rect 53228 51326 53230 51378
rect 53282 51326 53566 51378
rect 53618 51326 53620 51378
rect 53228 51324 53620 51326
rect 53228 51314 53284 51324
rect 53564 51314 53620 51324
rect 52780 50766 52782 50818
rect 52834 50766 52836 50818
rect 52780 50754 52836 50766
rect 52892 50596 52948 50606
rect 52892 50502 52948 50540
rect 53900 50596 53956 51438
rect 58156 51490 58212 51502
rect 58156 51438 58158 51490
rect 58210 51438 58212 51490
rect 57932 51156 57988 51166
rect 57932 50818 57988 51100
rect 57932 50766 57934 50818
rect 57986 50766 57988 50818
rect 57932 50754 57988 50766
rect 53900 50530 53956 50540
rect 55580 50596 55636 50606
rect 55580 50502 55636 50540
rect 51884 50418 51940 50428
rect 52780 50484 52836 50494
rect 52780 50390 52836 50428
rect 58156 50484 58212 51438
rect 58156 50418 58212 50428
rect 58156 49924 58212 49934
rect 58156 49922 58324 49924
rect 58156 49870 58158 49922
rect 58210 49870 58324 49922
rect 58156 49868 58324 49870
rect 58156 49858 58212 49868
rect 58156 49138 58212 49150
rect 58156 49086 58158 49138
rect 58210 49086 58212 49138
rect 58156 48468 58212 49086
rect 58268 49140 58324 49868
rect 58268 49074 58324 49084
rect 58156 48402 58212 48412
rect 57932 47570 57988 47582
rect 57932 47518 57934 47570
rect 57986 47518 57988 47570
rect 53228 47460 53284 47470
rect 51100 46786 51268 46788
rect 51100 46734 51102 46786
rect 51154 46734 51268 46786
rect 51100 46732 51268 46734
rect 51324 47346 51380 47358
rect 51324 47294 51326 47346
rect 51378 47294 51380 47346
rect 51100 46722 51156 46732
rect 49868 46610 49924 46620
rect 50652 46676 50708 46686
rect 50652 46582 50708 46620
rect 51324 46676 51380 47294
rect 52444 46786 52500 46798
rect 52444 46734 52446 46786
rect 52498 46734 52500 46786
rect 51324 46582 51380 46620
rect 51436 46674 51492 46686
rect 51436 46622 51438 46674
rect 51490 46622 51492 46674
rect 48188 46564 48244 46574
rect 48188 46470 48244 46508
rect 49532 46564 49588 46574
rect 46844 46396 47124 46452
rect 46844 45892 46900 45902
rect 46732 45836 46844 45892
rect 46844 45798 46900 45836
rect 47068 45890 47124 46396
rect 47068 45838 47070 45890
rect 47122 45838 47124 45890
rect 47068 45826 47124 45838
rect 49532 45892 49588 46508
rect 49532 45890 49700 45892
rect 49532 45838 49534 45890
rect 49586 45838 49700 45890
rect 49532 45836 49700 45838
rect 49532 45826 49588 45836
rect 46732 45668 46788 45678
rect 46620 45666 46788 45668
rect 46620 45614 46734 45666
rect 46786 45614 46788 45666
rect 46620 45612 46788 45614
rect 46732 45602 46788 45612
rect 44996 45500 45220 45556
rect 44940 45490 44996 45500
rect 44828 45330 45108 45332
rect 44828 45278 44830 45330
rect 44882 45278 45108 45330
rect 44828 45276 45108 45278
rect 44828 45266 44884 45276
rect 44604 45108 44660 45118
rect 44268 45106 44660 45108
rect 44268 45054 44606 45106
rect 44658 45054 44660 45106
rect 44268 45052 44660 45054
rect 44604 43540 44660 45052
rect 44940 43540 44996 43550
rect 44604 43538 44996 43540
rect 44604 43486 44942 43538
rect 44994 43486 44996 43538
rect 44604 43484 44996 43486
rect 44940 42868 44996 43484
rect 44940 42802 44996 42812
rect 44828 42532 44884 42542
rect 44492 41748 44548 41758
rect 44492 41654 44548 41692
rect 44828 41298 44884 42476
rect 45052 42532 45108 45276
rect 46396 45218 46452 45230
rect 46396 45166 46398 45218
rect 46450 45166 46452 45218
rect 46284 45108 46340 45118
rect 46172 45106 46340 45108
rect 46172 45054 46286 45106
rect 46338 45054 46340 45106
rect 46172 45052 46340 45054
rect 46172 44548 46228 45052
rect 46284 45042 46340 45052
rect 46172 44434 46228 44492
rect 46172 44382 46174 44434
rect 46226 44382 46228 44434
rect 46172 44370 46228 44382
rect 45948 44324 46004 44334
rect 45948 44230 46004 44268
rect 46396 44324 46452 45166
rect 46620 45108 46676 45118
rect 49644 45108 49700 45836
rect 49868 45890 49924 45902
rect 49868 45838 49870 45890
rect 49922 45838 49924 45890
rect 49756 45108 49812 45118
rect 46620 45106 47012 45108
rect 46620 45054 46622 45106
rect 46674 45054 47012 45106
rect 46620 45052 47012 45054
rect 49644 45106 49812 45108
rect 49644 45054 49758 45106
rect 49810 45054 49812 45106
rect 49644 45052 49812 45054
rect 46620 45042 46676 45052
rect 46396 44258 46452 44268
rect 46844 44324 46900 44334
rect 46844 44230 46900 44268
rect 46956 43540 47012 45052
rect 49756 45042 49812 45052
rect 47404 44996 47460 45006
rect 47404 44322 47460 44940
rect 49532 44994 49588 45006
rect 49532 44942 49534 44994
rect 49586 44942 49588 44994
rect 49532 44884 49588 44942
rect 49868 44884 49924 45838
rect 50316 45892 50372 45902
rect 50316 45798 50372 45836
rect 51324 45780 51380 45790
rect 51436 45780 51492 46622
rect 51660 46564 51716 46574
rect 51660 46114 51716 46508
rect 51660 46062 51662 46114
rect 51714 46062 51716 46114
rect 51660 46050 51716 46062
rect 51660 45892 51716 45902
rect 51324 45778 51492 45780
rect 51324 45726 51326 45778
rect 51378 45726 51492 45778
rect 51324 45724 51492 45726
rect 51548 45836 51660 45892
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 51324 45332 51380 45724
rect 50428 45276 51380 45332
rect 49532 44828 49924 44884
rect 50092 44884 50148 44894
rect 47740 44772 47796 44782
rect 47404 44270 47406 44322
rect 47458 44270 47460 44322
rect 47404 43762 47460 44270
rect 47404 43710 47406 43762
rect 47458 43710 47460 43762
rect 47404 43698 47460 43710
rect 47516 44434 47572 44446
rect 47516 44382 47518 44434
rect 47570 44382 47572 44434
rect 47516 44324 47572 44382
rect 47516 43764 47572 44268
rect 47628 43764 47684 43774
rect 47516 43762 47684 43764
rect 47516 43710 47630 43762
rect 47682 43710 47684 43762
rect 47516 43708 47684 43710
rect 47628 43698 47684 43708
rect 47068 43540 47124 43550
rect 46956 43538 47124 43540
rect 46956 43486 47070 43538
rect 47122 43486 47124 43538
rect 46956 43484 47124 43486
rect 47068 43474 47124 43484
rect 47516 43540 47572 43550
rect 47740 43540 47796 44716
rect 49532 44772 49588 44828
rect 50092 44790 50148 44828
rect 49532 44706 49588 44716
rect 48300 44210 48356 44222
rect 48300 44158 48302 44210
rect 48354 44158 48356 44210
rect 48300 43652 48356 44158
rect 50428 43764 50484 45276
rect 51548 45220 51604 45836
rect 51660 45798 51716 45836
rect 52444 45892 52500 46734
rect 52444 45826 52500 45836
rect 52892 46674 52948 46686
rect 52892 46622 52894 46674
rect 52946 46622 52948 46674
rect 52892 45890 52948 46622
rect 53116 46564 53172 46574
rect 53116 46470 53172 46508
rect 52892 45838 52894 45890
rect 52946 45838 52948 45890
rect 52892 45826 52948 45838
rect 53116 45780 53172 45790
rect 53228 45780 53284 47404
rect 55580 47460 55636 47470
rect 55580 47366 55636 47404
rect 57932 47124 57988 47518
rect 57932 47058 57988 47068
rect 53340 46676 53396 46686
rect 53340 46582 53396 46620
rect 53116 45778 53284 45780
rect 53116 45726 53118 45778
rect 53170 45726 53284 45778
rect 53116 45724 53284 45726
rect 53116 45714 53172 45724
rect 51212 45164 51604 45220
rect 50876 44884 50932 44894
rect 50876 44546 50932 44828
rect 50876 44494 50878 44546
rect 50930 44494 50932 44546
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50540 43764 50596 43774
rect 50428 43762 50596 43764
rect 50428 43710 50542 43762
rect 50594 43710 50596 43762
rect 50428 43708 50596 43710
rect 50540 43698 50596 43708
rect 50876 43708 50932 44494
rect 51212 44322 51268 45164
rect 57932 44434 57988 44446
rect 57932 44382 57934 44434
rect 57986 44382 57988 44434
rect 51212 44270 51214 44322
rect 51266 44270 51268 44322
rect 51212 44258 51268 44270
rect 53004 44324 53060 44334
rect 52668 44210 52724 44222
rect 52668 44158 52670 44210
rect 52722 44158 52724 44210
rect 50988 44098 51044 44110
rect 50988 44046 50990 44098
rect 51042 44046 51044 44098
rect 50988 43876 51044 44046
rect 50988 43820 51156 43876
rect 49756 43652 49812 43662
rect 48300 43586 48356 43596
rect 49644 43596 49756 43652
rect 47516 43538 47796 43540
rect 47516 43486 47518 43538
rect 47570 43486 47796 43538
rect 47516 43484 47796 43486
rect 47516 43474 47572 43484
rect 45052 42466 45108 42476
rect 45164 43426 45220 43438
rect 45164 43374 45166 43426
rect 45218 43374 45220 43426
rect 44828 41246 44830 41298
rect 44882 41246 44884 41298
rect 44828 41234 44884 41246
rect 45164 41300 45220 43374
rect 45276 43316 45332 43326
rect 45276 42756 45332 43260
rect 49532 43314 49588 43326
rect 49532 43262 49534 43314
rect 49586 43262 49588 43314
rect 45388 42756 45444 42766
rect 45276 42754 45444 42756
rect 45276 42702 45390 42754
rect 45442 42702 45444 42754
rect 45276 42700 45444 42702
rect 45276 42532 45332 42542
rect 45276 42196 45332 42476
rect 45388 42308 45444 42700
rect 45500 42756 45556 42766
rect 46172 42756 46228 42766
rect 49196 42756 49252 42766
rect 49532 42756 49588 43262
rect 45500 42754 46228 42756
rect 45500 42702 45502 42754
rect 45554 42702 46174 42754
rect 46226 42702 46228 42754
rect 45500 42700 46228 42702
rect 45500 42690 45556 42700
rect 46172 42690 46228 42700
rect 46732 42700 47012 42756
rect 46732 42642 46788 42700
rect 46732 42590 46734 42642
rect 46786 42590 46788 42642
rect 46732 42578 46788 42590
rect 45612 42532 45668 42542
rect 45612 42438 45668 42476
rect 45836 42530 45892 42542
rect 46508 42532 46564 42542
rect 45836 42478 45838 42530
rect 45890 42478 45892 42530
rect 45388 42252 45668 42308
rect 45276 42140 45444 42196
rect 45388 41970 45444 42140
rect 45388 41918 45390 41970
rect 45442 41918 45444 41970
rect 45388 41906 45444 41918
rect 45612 41970 45668 42252
rect 45612 41918 45614 41970
rect 45666 41918 45668 41970
rect 45612 41906 45668 41918
rect 45836 41748 45892 42478
rect 46284 42530 46676 42532
rect 46284 42478 46510 42530
rect 46562 42478 46676 42530
rect 46284 42476 46676 42478
rect 46284 42194 46340 42476
rect 46508 42466 46564 42476
rect 46284 42142 46286 42194
rect 46338 42142 46340 42194
rect 46284 42130 46340 42142
rect 46620 42084 46676 42476
rect 46844 42530 46900 42542
rect 46844 42478 46846 42530
rect 46898 42478 46900 42530
rect 46620 42028 46788 42084
rect 46620 41860 46676 41870
rect 45836 41654 45892 41692
rect 45948 41858 46676 41860
rect 45948 41806 46622 41858
rect 46674 41806 46676 41858
rect 45948 41804 46676 41806
rect 45948 41524 46004 41804
rect 46620 41794 46676 41804
rect 46732 41748 46788 42028
rect 46844 41972 46900 42478
rect 46844 41906 46900 41916
rect 46844 41748 46900 41758
rect 46732 41746 46900 41748
rect 46732 41694 46846 41746
rect 46898 41694 46900 41746
rect 46732 41692 46900 41694
rect 46844 41682 46900 41692
rect 45388 41468 46004 41524
rect 45388 41410 45444 41468
rect 46956 41412 47012 42700
rect 49196 42754 49588 42756
rect 49196 42702 49198 42754
rect 49250 42702 49588 42754
rect 49196 42700 49588 42702
rect 49644 42754 49700 43596
rect 49756 43558 49812 43596
rect 50652 43652 50708 43662
rect 50876 43652 51044 43708
rect 50652 43650 50820 43652
rect 50652 43598 50654 43650
rect 50706 43598 50820 43650
rect 50652 43596 50820 43598
rect 50652 43586 50708 43596
rect 50428 43538 50484 43550
rect 50428 43486 50430 43538
rect 50482 43486 50484 43538
rect 49868 43316 49924 43326
rect 49868 43222 49924 43260
rect 49644 42702 49646 42754
rect 49698 42702 49700 42754
rect 47180 42196 47236 42206
rect 47180 42102 47236 42140
rect 49196 42196 49252 42700
rect 49644 42690 49700 42702
rect 50092 42756 50148 42766
rect 50092 42662 50148 42700
rect 50428 42642 50484 43486
rect 50428 42590 50430 42642
rect 50482 42590 50484 42642
rect 50428 42532 50484 42590
rect 49196 42130 49252 42140
rect 50316 42476 50484 42532
rect 50652 43428 50708 43438
rect 50652 42530 50708 43372
rect 50652 42478 50654 42530
rect 50706 42478 50708 42530
rect 48412 41972 48468 41982
rect 45388 41358 45390 41410
rect 45442 41358 45444 41410
rect 45388 41346 45444 41358
rect 46396 41356 47012 41412
rect 47404 41748 47460 41758
rect 45164 41234 45220 41244
rect 45948 41300 46004 41310
rect 45948 41206 46004 41244
rect 45052 41186 45108 41198
rect 45052 41134 45054 41186
rect 45106 41134 45108 41186
rect 45052 40292 45108 41134
rect 46396 41076 46452 41356
rect 47404 41186 47460 41692
rect 47404 41134 47406 41186
rect 47458 41134 47460 41186
rect 47404 41122 47460 41134
rect 48412 41186 48468 41916
rect 50204 41860 50260 41870
rect 50316 41860 50372 42476
rect 50652 42466 50708 42478
rect 50764 42756 50820 43596
rect 50988 43426 51044 43652
rect 51100 43540 51156 43820
rect 51100 43474 51156 43484
rect 51212 43538 51268 43550
rect 51212 43486 51214 43538
rect 51266 43486 51268 43538
rect 50988 43374 50990 43426
rect 51042 43374 51044 43426
rect 50988 43362 51044 43374
rect 50764 42532 50820 42700
rect 50876 43316 50932 43326
rect 50876 42754 50932 43260
rect 51212 43316 51268 43486
rect 52332 43540 52388 43550
rect 52332 43446 52388 43484
rect 52444 43428 52500 43438
rect 52444 43334 52500 43372
rect 51212 43250 51268 43260
rect 52668 43314 52724 44158
rect 53004 44210 53060 44268
rect 55580 44324 55636 44334
rect 55580 44230 55636 44268
rect 53004 44158 53006 44210
rect 53058 44158 53060 44210
rect 53004 44146 53060 44158
rect 57932 43764 57988 44382
rect 57932 43698 57988 43708
rect 52668 43262 52670 43314
rect 52722 43262 52724 43314
rect 52668 43250 52724 43262
rect 57932 42866 57988 42878
rect 57932 42814 57934 42866
rect 57986 42814 57988 42866
rect 50876 42702 50878 42754
rect 50930 42702 50932 42754
rect 50876 42690 50932 42702
rect 51772 42756 51828 42766
rect 50764 42476 50932 42532
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50876 42196 50932 42476
rect 50652 42140 50932 42196
rect 51772 42194 51828 42700
rect 55580 42756 55636 42766
rect 55580 42662 55636 42700
rect 51772 42142 51774 42194
rect 51826 42142 51828 42194
rect 50652 41970 50708 42140
rect 51772 42130 51828 42142
rect 50652 41918 50654 41970
rect 50706 41918 50708 41970
rect 50652 41906 50708 41918
rect 51100 41972 51156 41982
rect 51436 41972 51492 41982
rect 51100 41970 51492 41972
rect 51100 41918 51102 41970
rect 51154 41918 51438 41970
rect 51490 41918 51492 41970
rect 51100 41916 51492 41918
rect 51100 41906 51156 41916
rect 51436 41906 51492 41916
rect 50204 41858 50372 41860
rect 50204 41806 50206 41858
rect 50258 41806 50372 41858
rect 50204 41804 50372 41806
rect 49532 41298 49588 41310
rect 49532 41246 49534 41298
rect 49586 41246 49588 41298
rect 48412 41134 48414 41186
rect 48466 41134 48468 41186
rect 48412 41122 48468 41134
rect 49196 41186 49252 41198
rect 49196 41134 49198 41186
rect 49250 41134 49252 41186
rect 45052 40226 45108 40236
rect 45724 41074 46452 41076
rect 45724 41022 46398 41074
rect 46450 41022 46452 41074
rect 45724 41020 46452 41022
rect 45724 39842 45780 41020
rect 46396 41010 46452 41020
rect 48076 41074 48132 41086
rect 48076 41022 48078 41074
rect 48130 41022 48132 41074
rect 48076 40964 48132 41022
rect 48076 40898 48132 40908
rect 45724 39790 45726 39842
rect 45778 39790 45780 39842
rect 45724 39778 45780 39790
rect 47852 40404 47908 40414
rect 45388 39620 45444 39630
rect 45388 39526 45444 39564
rect 46284 39620 46340 39630
rect 45164 39508 45220 39518
rect 45164 39414 45220 39452
rect 46284 39060 46340 39564
rect 46396 39618 46452 39630
rect 46396 39566 46398 39618
rect 46450 39566 46452 39618
rect 46396 39172 46452 39566
rect 46620 39620 46676 39630
rect 46620 39526 46676 39564
rect 46844 39620 46900 39630
rect 46844 39618 47012 39620
rect 46844 39566 46846 39618
rect 46898 39566 47012 39618
rect 46844 39564 47012 39566
rect 46844 39554 46900 39564
rect 46508 39396 46564 39406
rect 46508 39394 46900 39396
rect 46508 39342 46510 39394
rect 46562 39342 46900 39394
rect 46508 39340 46900 39342
rect 46508 39330 46564 39340
rect 46396 39116 46564 39172
rect 46284 38966 46340 39004
rect 44268 38836 44324 38846
rect 44268 36484 44324 38780
rect 45836 38834 45892 38846
rect 45836 38782 45838 38834
rect 45890 38782 45892 38834
rect 45836 37492 45892 38782
rect 46396 38836 46452 38846
rect 46396 38742 46452 38780
rect 46508 38834 46564 39116
rect 46508 38782 46510 38834
rect 46562 38782 46564 38834
rect 46508 38724 46564 38782
rect 46732 39060 46788 39070
rect 46508 38612 46676 38668
rect 45836 37426 45892 37436
rect 44380 37266 44436 37278
rect 44380 37214 44382 37266
rect 44434 37214 44436 37266
rect 44380 36706 44436 37214
rect 46620 37156 46676 38612
rect 46732 37378 46788 39004
rect 46844 38834 46900 39340
rect 46844 38782 46846 38834
rect 46898 38782 46900 38834
rect 46844 38770 46900 38782
rect 46956 38668 47012 39564
rect 47516 38946 47572 38958
rect 47516 38894 47518 38946
rect 47570 38894 47572 38946
rect 47404 38836 47460 38846
rect 47404 38742 47460 38780
rect 47516 38668 47572 38894
rect 46844 38612 47012 38668
rect 47180 38612 47572 38668
rect 47852 38722 47908 40348
rect 49084 40404 49140 40414
rect 49196 40404 49252 41134
rect 49140 40348 49252 40404
rect 49532 40964 49588 41246
rect 49868 41076 49924 41086
rect 50204 41076 50260 41804
rect 57932 41748 57988 42814
rect 57932 41682 57988 41692
rect 57932 41298 57988 41310
rect 57932 41246 57934 41298
rect 57986 41246 57988 41298
rect 49868 41074 50260 41076
rect 49868 41022 49870 41074
rect 49922 41022 50260 41074
rect 49868 41020 50260 41022
rect 50428 41188 50484 41198
rect 49868 41010 49924 41020
rect 49532 40402 49588 40908
rect 50428 40626 50484 41132
rect 55580 41188 55636 41198
rect 55580 41094 55636 41132
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50428 40574 50430 40626
rect 50482 40574 50484 40626
rect 50428 40562 50484 40574
rect 49532 40350 49534 40402
rect 49586 40350 49588 40402
rect 49084 40310 49140 40348
rect 49532 40338 49588 40350
rect 49756 40404 49812 40414
rect 50092 40404 50148 40414
rect 49756 40402 50148 40404
rect 49756 40350 49758 40402
rect 49810 40350 50094 40402
rect 50146 40350 50148 40402
rect 49756 40348 50148 40350
rect 49756 40338 49812 40348
rect 50092 40338 50148 40348
rect 57932 40404 57988 41246
rect 57932 40338 57988 40348
rect 58156 39396 58212 39406
rect 58156 39394 58324 39396
rect 58156 39342 58158 39394
rect 58210 39342 58324 39394
rect 58156 39340 58324 39342
rect 58156 39330 58212 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 58268 39060 58324 39340
rect 58268 38994 58324 39004
rect 47852 38670 47854 38722
rect 47906 38670 47908 38722
rect 47852 38658 47908 38670
rect 58156 38946 58212 38958
rect 58156 38894 58158 38946
rect 58210 38894 58212 38946
rect 46844 38162 46900 38612
rect 46844 38110 46846 38162
rect 46898 38110 46900 38162
rect 46844 37492 46900 38110
rect 46844 37426 46900 37436
rect 47180 37938 47236 38612
rect 58156 38388 58212 38894
rect 58156 38322 58212 38332
rect 57932 38162 57988 38174
rect 57932 38110 57934 38162
rect 57986 38110 57988 38162
rect 48188 38052 48244 38062
rect 47180 37886 47182 37938
rect 47234 37886 47236 37938
rect 46732 37326 46734 37378
rect 46786 37326 46788 37378
rect 46732 37314 46788 37326
rect 46956 37156 47012 37166
rect 46620 37154 47012 37156
rect 46620 37102 46958 37154
rect 47010 37102 47012 37154
rect 46620 37100 47012 37102
rect 46956 37090 47012 37100
rect 44380 36654 44382 36706
rect 44434 36654 44436 36706
rect 44380 36642 44436 36654
rect 47180 36708 47236 37886
rect 47404 38050 48244 38052
rect 47404 37998 48190 38050
rect 48242 37998 48244 38050
rect 47404 37996 48244 37998
rect 47292 37492 47348 37502
rect 47404 37492 47460 37996
rect 48188 37986 48244 37996
rect 49532 38052 49588 38062
rect 48860 37940 48916 37950
rect 49196 37940 49252 37950
rect 48860 37938 49252 37940
rect 48860 37886 48862 37938
rect 48914 37886 49198 37938
rect 49250 37886 49252 37938
rect 48860 37884 49252 37886
rect 48860 37874 48916 37884
rect 49196 37874 49252 37884
rect 49532 37938 49588 37996
rect 55580 38052 55636 38062
rect 55580 37958 55636 37996
rect 49532 37886 49534 37938
rect 49586 37886 49588 37938
rect 49532 37874 49588 37886
rect 57932 37716 57988 38110
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 57932 37650 57988 37660
rect 50556 37594 50820 37604
rect 47292 37490 47460 37492
rect 47292 37438 47294 37490
rect 47346 37438 47460 37490
rect 47292 37436 47460 37438
rect 47292 37426 47348 37436
rect 47404 36708 47460 36718
rect 47180 36706 47460 36708
rect 47180 36654 47406 36706
rect 47458 36654 47460 36706
rect 47180 36652 47460 36654
rect 47404 36642 47460 36652
rect 45612 36596 45668 36606
rect 45612 36502 45668 36540
rect 47068 36596 47124 36606
rect 47068 36502 47124 36540
rect 57932 36594 57988 36606
rect 57932 36542 57934 36594
rect 57986 36542 57988 36594
rect 44268 36428 44436 36484
rect 44268 36260 44324 36270
rect 44212 36258 44324 36260
rect 44212 36206 44270 36258
rect 44322 36206 44324 36258
rect 44212 36204 44324 36206
rect 44156 36166 44212 36204
rect 44268 36194 44324 36204
rect 43932 35646 43934 35698
rect 43986 35646 43988 35698
rect 43932 35634 43988 35646
rect 43372 34302 43374 34354
rect 43426 34302 43428 34354
rect 43372 34290 43428 34302
rect 44156 35028 44212 35038
rect 43148 34130 43204 34142
rect 43148 34078 43150 34130
rect 43202 34078 43204 34130
rect 42140 33294 42142 33346
rect 42194 33294 42196 33346
rect 42140 33236 42196 33294
rect 42140 33170 42196 33180
rect 42252 33292 42980 33348
rect 38892 32956 39508 33012
rect 38892 32900 38948 32956
rect 38668 32722 38724 32732
rect 38780 32844 38948 32900
rect 38780 32562 38836 32844
rect 39004 32788 39060 32798
rect 39004 32676 39060 32732
rect 39452 32786 39508 32956
rect 41916 33122 41972 33134
rect 41916 33070 41918 33122
rect 41970 33070 41972 33122
rect 39452 32734 39454 32786
rect 39506 32734 39508 32786
rect 39452 32722 39508 32734
rect 39676 32788 39732 32798
rect 39676 32786 40180 32788
rect 39676 32734 39678 32786
rect 39730 32734 40180 32786
rect 39676 32732 40180 32734
rect 39676 32722 39732 32732
rect 39116 32676 39172 32686
rect 39004 32674 39172 32676
rect 39004 32622 39118 32674
rect 39170 32622 39172 32674
rect 39004 32620 39172 32622
rect 39116 32610 39172 32620
rect 38780 32510 38782 32562
rect 38834 32510 38836 32562
rect 38780 32498 38836 32510
rect 38892 32562 38948 32574
rect 38892 32510 38894 32562
rect 38946 32510 38948 32562
rect 38892 32452 38948 32510
rect 39228 32564 39284 32574
rect 39228 32470 39284 32508
rect 39676 32564 39732 32574
rect 39788 32564 39844 32574
rect 39732 32562 39844 32564
rect 39732 32510 39790 32562
rect 39842 32510 39844 32562
rect 39732 32508 39844 32510
rect 38892 32386 38948 32396
rect 38556 32060 38836 32116
rect 37100 31892 37380 31948
rect 37660 31892 38276 31948
rect 36988 30258 37044 30268
rect 35868 30046 35870 30098
rect 35922 30046 35924 30098
rect 35868 30034 35924 30046
rect 35868 29764 35924 29774
rect 35756 29708 35868 29764
rect 33516 28644 33572 28654
rect 34076 28644 34132 28654
rect 33516 28642 34132 28644
rect 33516 28590 33518 28642
rect 33570 28590 34078 28642
rect 34130 28590 34132 28642
rect 33516 28588 34132 28590
rect 33516 28578 33572 28588
rect 34076 28578 34132 28588
rect 34412 28644 34468 29596
rect 34412 28578 34468 28588
rect 34972 29426 35028 29438
rect 34972 29374 34974 29426
rect 35026 29374 35028 29426
rect 33740 28420 33796 28430
rect 33740 28418 34132 28420
rect 33740 28366 33742 28418
rect 33794 28366 34132 28418
rect 33740 28364 34132 28366
rect 33740 28354 33796 28364
rect 33068 27468 33236 27524
rect 31724 26338 31780 26348
rect 30828 26292 30884 26302
rect 29036 26180 29092 26190
rect 29036 26086 29092 26124
rect 29708 25732 29764 25742
rect 29708 25638 29764 25676
rect 30380 25732 30436 25742
rect 28308 25452 28532 25508
rect 29484 25508 29540 25518
rect 27580 25394 27636 25406
rect 27580 25342 27582 25394
rect 27634 25342 27636 25394
rect 27580 25284 27636 25342
rect 28252 25394 28308 25452
rect 29484 25414 29540 25452
rect 29932 25508 29988 25518
rect 30380 25508 30436 25676
rect 30828 25620 30884 26236
rect 29932 25506 30436 25508
rect 29932 25454 29934 25506
rect 29986 25454 30382 25506
rect 30434 25454 30436 25506
rect 29932 25452 30436 25454
rect 29932 25442 29988 25452
rect 30380 25442 30436 25452
rect 30716 25618 30884 25620
rect 30716 25566 30830 25618
rect 30882 25566 30884 25618
rect 30716 25564 30884 25566
rect 30716 25508 30772 25564
rect 30828 25554 30884 25564
rect 31052 26178 31108 26190
rect 31052 26126 31054 26178
rect 31106 26126 31108 26178
rect 31052 25508 31108 26126
rect 31276 25508 31332 25518
rect 31052 25506 31332 25508
rect 31052 25454 31278 25506
rect 31330 25454 31332 25506
rect 31052 25452 31332 25454
rect 28252 25342 28254 25394
rect 28306 25342 28308 25394
rect 28252 25330 28308 25342
rect 27244 25282 27636 25284
rect 27244 25230 27246 25282
rect 27298 25230 27636 25282
rect 27244 25228 27636 25230
rect 27692 25284 27748 25294
rect 28588 25284 28644 25294
rect 26684 23762 26740 23772
rect 26908 24722 26964 24734
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26908 23380 26964 24670
rect 27132 23940 27188 23950
rect 27132 23846 27188 23884
rect 27244 23548 27300 25228
rect 27692 25190 27748 25228
rect 28476 25282 28644 25284
rect 28476 25230 28590 25282
rect 28642 25230 28644 25282
rect 28476 25228 28644 25230
rect 28028 24724 28084 24734
rect 27580 23828 27636 23838
rect 27580 23734 27636 23772
rect 28028 23826 28084 24668
rect 28140 24722 28196 24734
rect 28476 24724 28532 25228
rect 28588 25218 28644 25228
rect 28700 25284 28756 25294
rect 28140 24670 28142 24722
rect 28194 24670 28196 24722
rect 28140 24276 28196 24670
rect 28140 24210 28196 24220
rect 28252 24722 28532 24724
rect 28252 24670 28478 24722
rect 28530 24670 28532 24722
rect 28252 24668 28532 24670
rect 28028 23774 28030 23826
rect 28082 23774 28084 23826
rect 26908 23286 26964 23324
rect 27132 23492 27300 23548
rect 26684 23154 26740 23166
rect 26684 23102 26686 23154
rect 26738 23102 26740 23154
rect 26684 23044 26740 23102
rect 27020 23156 27076 23166
rect 27020 23062 27076 23100
rect 26684 22978 26740 22988
rect 27132 22484 27188 23492
rect 27468 23268 27524 23278
rect 27468 23154 27524 23212
rect 27468 23102 27470 23154
rect 27522 23102 27524 23154
rect 27468 23090 27524 23102
rect 27692 23156 27748 23166
rect 28028 23156 28084 23774
rect 28140 23938 28196 23950
rect 28140 23886 28142 23938
rect 28194 23886 28196 23938
rect 28140 23380 28196 23886
rect 28140 23314 28196 23324
rect 28028 23100 28196 23156
rect 27692 23062 27748 23100
rect 28028 22932 28084 22942
rect 28028 22838 28084 22876
rect 26572 22306 26628 22316
rect 26908 22428 27188 22484
rect 27804 22484 27860 22522
rect 26684 21698 26740 21710
rect 26684 21646 26686 21698
rect 26738 21646 26740 21698
rect 26572 21474 26628 21486
rect 26572 21422 26574 21474
rect 26626 21422 26628 21474
rect 26572 20804 26628 21422
rect 26572 20738 26628 20748
rect 26572 20580 26628 20590
rect 26572 20486 26628 20524
rect 26460 20300 26628 20356
rect 26236 20018 26404 20020
rect 26236 19966 26238 20018
rect 26290 19966 26404 20018
rect 26236 19964 26404 19966
rect 26236 19954 26292 19964
rect 26348 18788 26404 19964
rect 26460 19236 26516 19246
rect 26460 19142 26516 19180
rect 26348 18722 26404 18732
rect 26124 18620 26292 18676
rect 25788 18610 25844 18620
rect 25676 18510 25678 18562
rect 25730 18510 25732 18562
rect 25676 18498 25732 18510
rect 25900 18564 25956 18574
rect 25564 18386 25620 18396
rect 25340 17836 25844 17892
rect 25172 17612 25620 17668
rect 25116 17574 25172 17612
rect 25228 17442 25284 17454
rect 25452 17444 25508 17454
rect 25228 17390 25230 17442
rect 25282 17390 25284 17442
rect 25228 17220 25284 17390
rect 25228 17154 25284 17164
rect 25340 17442 25508 17444
rect 25340 17390 25454 17442
rect 25506 17390 25508 17442
rect 25340 17388 25508 17390
rect 25004 16548 25060 16558
rect 25004 16098 25060 16492
rect 25340 16324 25396 17388
rect 25452 17378 25508 17388
rect 25564 16882 25620 17612
rect 25564 16830 25566 16882
rect 25618 16830 25620 16882
rect 25564 16818 25620 16830
rect 25676 16884 25732 16894
rect 25676 16770 25732 16828
rect 25676 16718 25678 16770
rect 25730 16718 25732 16770
rect 25676 16706 25732 16718
rect 25676 16436 25732 16446
rect 25340 16268 25620 16324
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 25004 16034 25060 16046
rect 25340 16100 25396 16110
rect 25340 15540 25396 16044
rect 25228 15538 25396 15540
rect 25228 15486 25342 15538
rect 25394 15486 25396 15538
rect 25228 15484 25396 15486
rect 24892 15092 25060 15148
rect 24892 14420 24948 14430
rect 24892 14326 24948 14364
rect 25004 14196 25060 15092
rect 24724 13916 24836 13972
rect 24892 14140 25060 14196
rect 24668 13878 24724 13916
rect 24780 12852 24836 12862
rect 24556 12850 24836 12852
rect 24556 12798 24782 12850
rect 24834 12798 24836 12850
rect 24556 12796 24836 12798
rect 24780 12786 24836 12796
rect 24556 12178 24612 12190
rect 24556 12126 24558 12178
rect 24610 12126 24612 12178
rect 24108 11900 24388 11956
rect 24220 11396 24276 11406
rect 24108 10836 24164 10846
rect 24108 9492 24164 10780
rect 24220 10834 24276 11340
rect 24332 11394 24388 11900
rect 24444 11954 24500 11966
rect 24444 11902 24446 11954
rect 24498 11902 24500 11954
rect 24444 11506 24500 11902
rect 24444 11454 24446 11506
rect 24498 11454 24500 11506
rect 24444 11442 24500 11454
rect 24332 11342 24334 11394
rect 24386 11342 24388 11394
rect 24332 11330 24388 11342
rect 24220 10782 24222 10834
rect 24274 10782 24276 10834
rect 24220 10770 24276 10782
rect 24556 10836 24612 12126
rect 24892 10836 24948 14140
rect 25228 13524 25284 15484
rect 25340 15474 25396 15484
rect 25564 15148 25620 16268
rect 25676 15876 25732 16380
rect 25788 16100 25844 17836
rect 25900 16994 25956 18508
rect 26124 18452 26180 18462
rect 25900 16942 25902 16994
rect 25954 16942 25956 16994
rect 25900 16930 25956 16942
rect 26012 18450 26180 18452
rect 26012 18398 26126 18450
rect 26178 18398 26180 18450
rect 26012 18396 26180 18398
rect 25788 16034 25844 16044
rect 25676 15820 25844 15876
rect 25676 15652 25732 15662
rect 25676 15314 25732 15596
rect 25788 15426 25844 15820
rect 25788 15374 25790 15426
rect 25842 15374 25844 15426
rect 25788 15362 25844 15374
rect 25676 15262 25678 15314
rect 25730 15262 25732 15314
rect 25676 15250 25732 15262
rect 25116 13412 25172 13422
rect 25004 13076 25060 13086
rect 25004 12962 25060 13020
rect 25116 13074 25172 13356
rect 25116 13022 25118 13074
rect 25170 13022 25172 13074
rect 25116 13010 25172 13022
rect 25004 12910 25006 12962
rect 25058 12910 25060 12962
rect 25004 11844 25060 12910
rect 25228 12740 25284 13468
rect 25340 15092 25620 15148
rect 25788 15204 25844 15214
rect 26012 15148 26068 18396
rect 26124 18386 26180 18396
rect 26236 17892 26292 18620
rect 26236 17836 26516 17892
rect 26236 17668 26292 17678
rect 26124 17442 26180 17454
rect 26124 17390 26126 17442
rect 26178 17390 26180 17442
rect 26124 17108 26180 17390
rect 26124 15316 26180 17052
rect 26236 16098 26292 17612
rect 26236 16046 26238 16098
rect 26290 16046 26292 16098
rect 26236 16034 26292 16046
rect 26348 16882 26404 16894
rect 26348 16830 26350 16882
rect 26402 16830 26404 16882
rect 26348 15538 26404 16830
rect 26460 16772 26516 17836
rect 26572 17442 26628 20300
rect 26684 20020 26740 21646
rect 26684 19954 26740 19964
rect 26796 19906 26852 19918
rect 26796 19854 26798 19906
rect 26850 19854 26852 19906
rect 26796 19460 26852 19854
rect 26796 19394 26852 19404
rect 26684 19236 26740 19246
rect 26684 19142 26740 19180
rect 26796 19234 26852 19246
rect 26796 19182 26798 19234
rect 26850 19182 26852 19234
rect 26796 18452 26852 19182
rect 26908 18564 26964 22428
rect 27804 22418 27860 22428
rect 27468 22372 27524 22382
rect 27468 22370 27636 22372
rect 27468 22318 27470 22370
rect 27522 22318 27636 22370
rect 27468 22316 27636 22318
rect 27468 22306 27524 22316
rect 27132 22260 27188 22298
rect 27188 22204 27412 22260
rect 27132 22194 27188 22204
rect 27132 22036 27188 22046
rect 27132 21700 27188 21980
rect 27356 21924 27412 22204
rect 27356 21868 27524 21924
rect 27468 21810 27524 21868
rect 27468 21758 27470 21810
rect 27522 21758 27524 21810
rect 27468 21746 27524 21758
rect 27356 21700 27412 21710
rect 27020 21698 27412 21700
rect 27020 21646 27358 21698
rect 27410 21646 27412 21698
rect 27020 21644 27412 21646
rect 27020 20914 27076 21644
rect 27356 21634 27412 21644
rect 27580 21588 27636 22316
rect 27804 22258 27860 22270
rect 27804 22206 27806 22258
rect 27858 22206 27860 22258
rect 27804 21924 27860 22206
rect 27804 21858 27860 21868
rect 27692 21812 27748 21822
rect 27692 21718 27748 21756
rect 27580 21532 27860 21588
rect 27580 21364 27636 21374
rect 27020 20862 27022 20914
rect 27074 20862 27076 20914
rect 27020 20850 27076 20862
rect 27244 20916 27300 20926
rect 27132 20132 27188 20142
rect 27244 20132 27300 20860
rect 27356 20580 27412 20590
rect 27356 20486 27412 20524
rect 27580 20242 27636 21308
rect 27580 20190 27582 20242
rect 27634 20190 27636 20242
rect 27580 20178 27636 20190
rect 27132 20130 27524 20132
rect 27132 20078 27134 20130
rect 27186 20078 27524 20130
rect 27132 20076 27524 20078
rect 27132 20066 27188 20076
rect 27356 19796 27412 19806
rect 27244 19794 27412 19796
rect 27244 19742 27358 19794
rect 27410 19742 27412 19794
rect 27244 19740 27412 19742
rect 27132 19124 27188 19134
rect 27132 19030 27188 19068
rect 26908 18508 27076 18564
rect 26796 18386 26852 18396
rect 26908 18338 26964 18350
rect 26908 18286 26910 18338
rect 26962 18286 26964 18338
rect 26908 18228 26964 18286
rect 26908 18162 26964 18172
rect 27020 17780 27076 18508
rect 27020 17778 27188 17780
rect 27020 17726 27022 17778
rect 27074 17726 27188 17778
rect 27020 17724 27188 17726
rect 27020 17714 27076 17724
rect 26572 17390 26574 17442
rect 26626 17390 26628 17442
rect 26572 16884 26628 17390
rect 26908 17444 26964 17454
rect 26908 17108 26964 17388
rect 27132 17220 27188 17724
rect 27244 17668 27300 19740
rect 27356 19730 27412 19740
rect 27244 17602 27300 17612
rect 27356 19572 27412 19582
rect 27356 17444 27412 19516
rect 27468 19346 27524 20076
rect 27468 19294 27470 19346
rect 27522 19294 27524 19346
rect 27468 19282 27524 19294
rect 27692 19234 27748 19246
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 19124 27748 19182
rect 27692 19058 27748 19068
rect 27692 18676 27748 18686
rect 27804 18676 27860 21532
rect 28028 21476 28084 21486
rect 27916 21474 28084 21476
rect 27916 21422 28030 21474
rect 28082 21422 28084 21474
rect 27916 21420 28084 21422
rect 27916 21140 27972 21420
rect 28028 21410 28084 21420
rect 28140 21252 28196 23100
rect 28252 22708 28308 24668
rect 28476 24658 28532 24668
rect 28700 24610 28756 25228
rect 29036 25284 29092 25294
rect 29036 25282 29876 25284
rect 29036 25230 29038 25282
rect 29090 25230 29876 25282
rect 29036 25228 29876 25230
rect 29036 25218 29092 25228
rect 29820 24834 29876 25228
rect 29820 24782 29822 24834
rect 29874 24782 29876 24834
rect 29820 24770 29876 24782
rect 30716 24722 30772 25452
rect 30716 24670 30718 24722
rect 30770 24670 30772 24722
rect 30716 24658 30772 24670
rect 30828 24724 30884 24734
rect 30828 24630 30884 24668
rect 31164 24724 31220 24734
rect 31276 24724 31332 25452
rect 31500 25508 31556 25518
rect 32844 25508 32900 25518
rect 31556 25452 31780 25508
rect 31500 25414 31556 25452
rect 31724 25172 31780 25452
rect 32844 25414 32900 25452
rect 32060 25394 32116 25406
rect 32060 25342 32062 25394
rect 32114 25342 32116 25394
rect 32060 25284 32116 25342
rect 32060 25218 32116 25228
rect 31724 25116 31892 25172
rect 31164 24722 31276 24724
rect 31164 24670 31166 24722
rect 31218 24670 31276 24722
rect 31164 24668 31276 24670
rect 28700 24558 28702 24610
rect 28754 24558 28756 24610
rect 28700 24546 28756 24558
rect 31052 24610 31108 24622
rect 31052 24558 31054 24610
rect 31106 24558 31108 24610
rect 28476 24498 28532 24510
rect 28476 24446 28478 24498
rect 28530 24446 28532 24498
rect 28364 24050 28420 24062
rect 28364 23998 28366 24050
rect 28418 23998 28420 24050
rect 28364 23492 28420 23998
rect 28364 23426 28420 23436
rect 28476 23268 28532 24446
rect 29932 24500 29988 24510
rect 29932 24498 30548 24500
rect 29932 24446 29934 24498
rect 29986 24446 30548 24498
rect 29932 24444 30548 24446
rect 29932 24434 29988 24444
rect 30044 24164 30100 24174
rect 30044 24050 30100 24108
rect 30044 23998 30046 24050
rect 30098 23998 30100 24050
rect 30044 23986 30100 23998
rect 30268 23940 30324 23950
rect 30268 23826 30324 23884
rect 30492 23938 30548 24444
rect 30492 23886 30494 23938
rect 30546 23886 30548 23938
rect 30492 23874 30548 23886
rect 30716 24164 30772 24174
rect 30268 23774 30270 23826
rect 30322 23774 30324 23826
rect 28364 23156 28420 23166
rect 28476 23156 28532 23212
rect 29484 23716 29540 23726
rect 28588 23156 28644 23166
rect 28476 23154 28644 23156
rect 28476 23102 28590 23154
rect 28642 23102 28644 23154
rect 28476 23100 28644 23102
rect 28364 23062 28420 23100
rect 28588 23090 28644 23100
rect 28252 22642 28308 22652
rect 28364 22820 28420 22830
rect 28252 22372 28308 22382
rect 28252 22278 28308 22316
rect 28364 21586 28420 22764
rect 29148 22260 29204 22270
rect 29148 21698 29204 22204
rect 29148 21646 29150 21698
rect 29202 21646 29204 21698
rect 29148 21634 29204 21646
rect 29372 22146 29428 22158
rect 29372 22094 29374 22146
rect 29426 22094 29428 22146
rect 28364 21534 28366 21586
rect 28418 21534 28420 21586
rect 28140 21196 28308 21252
rect 27916 21074 27972 21084
rect 28028 21028 28084 21038
rect 27916 20802 27972 20814
rect 27916 20750 27918 20802
rect 27970 20750 27972 20802
rect 27916 20468 27972 20750
rect 27916 20402 27972 20412
rect 28028 19236 28084 20972
rect 28140 19906 28196 19918
rect 28140 19854 28142 19906
rect 28194 19854 28196 19906
rect 28140 19460 28196 19854
rect 28252 19572 28308 21196
rect 28364 20580 28420 21534
rect 28364 20486 28420 20524
rect 28812 21586 28868 21598
rect 28812 21534 28814 21586
rect 28866 21534 28868 21586
rect 28812 20468 28868 21534
rect 29372 21588 29428 22094
rect 29372 21252 29428 21532
rect 29372 21186 29428 21196
rect 29372 20578 29428 20590
rect 29372 20526 29374 20578
rect 29426 20526 29428 20578
rect 29372 20468 29428 20526
rect 28476 19906 28532 19918
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28476 19794 28532 19854
rect 28476 19742 28478 19794
rect 28530 19742 28532 19794
rect 28476 19730 28532 19742
rect 28252 19516 28644 19572
rect 28196 19404 28532 19460
rect 28140 19394 28196 19404
rect 28476 19346 28532 19404
rect 28476 19294 28478 19346
rect 28530 19294 28532 19346
rect 28476 19282 28532 19294
rect 28028 19180 28308 19236
rect 28028 19012 28084 19022
rect 28028 18918 28084 18956
rect 27748 18620 27860 18676
rect 28140 18788 28196 18798
rect 27692 18562 27748 18620
rect 27692 18510 27694 18562
rect 27746 18510 27748 18562
rect 27580 18452 27636 18462
rect 27580 18358 27636 18396
rect 27356 17378 27412 17388
rect 27580 17442 27636 17454
rect 27580 17390 27582 17442
rect 27634 17390 27636 17442
rect 27132 17164 27524 17220
rect 26908 17106 27188 17108
rect 26908 17054 26910 17106
rect 26962 17054 27188 17106
rect 26908 17052 27188 17054
rect 26908 17042 26964 17052
rect 27132 16884 27188 17052
rect 26572 16828 27076 16884
rect 26460 15988 26516 16716
rect 26908 16324 26964 16334
rect 26572 16212 26628 16222
rect 26572 16118 26628 16156
rect 26460 15922 26516 15932
rect 26684 16100 26740 16110
rect 26348 15486 26350 15538
rect 26402 15486 26404 15538
rect 26348 15474 26404 15486
rect 26460 15652 26516 15662
rect 26684 15652 26740 16044
rect 26908 16098 26964 16268
rect 26908 16046 26910 16098
rect 26962 16046 26964 16098
rect 26908 16034 26964 16046
rect 26516 15596 26740 15652
rect 26124 15250 26180 15260
rect 26460 15148 26516 15596
rect 26796 15316 26852 15326
rect 27020 15316 27076 16828
rect 26796 15314 27076 15316
rect 26796 15262 26798 15314
rect 26850 15262 27076 15314
rect 26796 15260 27076 15262
rect 26796 15250 26852 15260
rect 25340 12852 25396 15092
rect 25788 14754 25844 15148
rect 25788 14702 25790 14754
rect 25842 14702 25844 14754
rect 25788 14690 25844 14702
rect 25900 15092 26068 15148
rect 26348 15092 26516 15148
rect 26572 15092 26628 15102
rect 25676 14532 25732 14542
rect 25452 14420 25508 14430
rect 25452 14418 25620 14420
rect 25452 14366 25454 14418
rect 25506 14366 25620 14418
rect 25452 14364 25620 14366
rect 25452 14354 25508 14364
rect 25452 13860 25508 13870
rect 25452 13766 25508 13804
rect 25564 13300 25620 14364
rect 25676 13970 25732 14476
rect 25676 13918 25678 13970
rect 25730 13918 25732 13970
rect 25676 13906 25732 13918
rect 25788 13860 25844 13870
rect 25788 13634 25844 13804
rect 25788 13582 25790 13634
rect 25842 13582 25844 13634
rect 25788 13570 25844 13582
rect 25900 13858 25956 15092
rect 26124 14642 26180 14654
rect 26124 14590 26126 14642
rect 26178 14590 26180 14642
rect 26012 14308 26068 14318
rect 26012 14214 26068 14252
rect 25900 13806 25902 13858
rect 25954 13806 25956 13858
rect 25564 13234 25620 13244
rect 25452 12852 25508 12862
rect 25340 12796 25452 12852
rect 25452 12786 25508 12796
rect 25228 12684 25396 12740
rect 25004 11732 25284 11788
rect 25116 11620 25172 11630
rect 25116 11526 25172 11564
rect 24892 10780 25060 10836
rect 24332 10610 24388 10622
rect 24332 10558 24334 10610
rect 24386 10558 24388 10610
rect 24108 9426 24164 9436
rect 24220 9828 24276 9838
rect 24108 9268 24164 9278
rect 23996 9266 24164 9268
rect 23996 9214 24110 9266
rect 24162 9214 24164 9266
rect 23996 9212 24164 9214
rect 24108 9202 24164 9212
rect 24220 9156 24276 9772
rect 24220 9090 24276 9100
rect 23884 8978 23940 8988
rect 24108 9042 24164 9054
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 23716 8652 23828 8708
rect 23660 8642 23716 8652
rect 23548 7534 23550 7586
rect 23602 7534 23604 7586
rect 23548 7522 23604 7534
rect 24108 7588 24164 8990
rect 23436 7310 23438 7362
rect 23490 7310 23492 7362
rect 23436 7298 23492 7310
rect 24108 6580 24164 7532
rect 24108 6514 24164 6524
rect 24220 8258 24276 8270
rect 24220 8206 24222 8258
rect 24274 8206 24276 8258
rect 24220 7364 24276 8206
rect 23436 6244 23492 6254
rect 23436 5682 23492 6188
rect 23436 5630 23438 5682
rect 23490 5630 23492 5682
rect 23436 5618 23492 5630
rect 24220 4676 24276 7308
rect 24332 8260 24388 10558
rect 24444 10164 24500 10174
rect 24556 10164 24612 10780
rect 25004 10724 25060 10780
rect 24668 10610 24724 10622
rect 24668 10558 24670 10610
rect 24722 10558 24724 10610
rect 24668 10500 24724 10558
rect 24668 10276 24724 10444
rect 24892 10612 24948 10622
rect 24668 10210 24724 10220
rect 24780 10388 24836 10398
rect 24500 10108 24612 10164
rect 24444 10098 24500 10108
rect 24668 10052 24724 10062
rect 24668 9938 24724 9996
rect 24668 9886 24670 9938
rect 24722 9886 24724 9938
rect 24668 9874 24724 9886
rect 24780 8484 24836 10332
rect 24668 8428 24836 8484
rect 24332 5572 24388 8204
rect 24556 8372 24612 8382
rect 24556 8146 24612 8316
rect 24556 8094 24558 8146
rect 24610 8094 24612 8146
rect 24556 8082 24612 8094
rect 24668 7812 24724 8428
rect 24556 7756 24724 7812
rect 24892 8370 24948 10556
rect 24892 8318 24894 8370
rect 24946 8318 24948 8370
rect 24444 7476 24500 7486
rect 24444 6916 24500 7420
rect 24556 7364 24612 7756
rect 24668 7588 24724 7598
rect 24892 7588 24948 8318
rect 24668 7586 24948 7588
rect 24668 7534 24670 7586
rect 24722 7534 24948 7586
rect 24668 7532 24948 7534
rect 24668 7522 24724 7532
rect 24556 7308 24836 7364
rect 24444 6850 24500 6860
rect 24668 6690 24724 6702
rect 24668 6638 24670 6690
rect 24722 6638 24724 6690
rect 24556 6132 24612 6142
rect 24556 6018 24612 6076
rect 24556 5966 24558 6018
rect 24610 5966 24612 6018
rect 24556 5954 24612 5966
rect 24332 5506 24388 5516
rect 24220 4610 24276 4620
rect 24332 5236 24388 5246
rect 23436 4338 23492 4350
rect 23436 4286 23438 4338
rect 23490 4286 23492 4338
rect 23436 4116 23492 4286
rect 23436 4050 23492 4060
rect 23996 4340 24052 4350
rect 23996 3666 24052 4284
rect 23996 3614 23998 3666
rect 24050 3614 24052 3666
rect 23996 3602 24052 3614
rect 23548 3556 23604 3566
rect 24332 3556 24388 5180
rect 24444 5122 24500 5134
rect 24444 5070 24446 5122
rect 24498 5070 24500 5122
rect 24444 5012 24500 5070
rect 24444 4946 24500 4956
rect 24556 3556 24612 3566
rect 24332 3554 24612 3556
rect 24332 3502 24558 3554
rect 24610 3502 24612 3554
rect 24332 3500 24612 3502
rect 23548 3462 23604 3500
rect 24556 3490 24612 3500
rect 23268 3388 23380 3444
rect 23212 3378 23268 3388
rect 22988 3332 23044 3342
rect 19516 2996 19572 3006
rect 19628 2996 19684 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20412 3108 20468 3332
rect 22876 3276 22988 3332
rect 22988 3266 23044 3276
rect 20412 3042 20468 3052
rect 19572 2940 19684 2996
rect 19516 2930 19572 2940
rect 18956 2706 19012 2716
rect 24668 2324 24724 6638
rect 24780 4562 24836 7308
rect 24892 5236 24948 5246
rect 25004 5236 25060 10668
rect 25228 10722 25284 11732
rect 25228 10670 25230 10722
rect 25282 10670 25284 10722
rect 25228 10658 25284 10670
rect 25116 9828 25172 9838
rect 25340 9828 25396 12684
rect 25676 11956 25732 11966
rect 25564 10724 25620 10734
rect 25116 9734 25172 9772
rect 25228 9772 25396 9828
rect 25452 10610 25508 10622
rect 25452 10558 25454 10610
rect 25506 10558 25508 10610
rect 25452 9940 25508 10558
rect 25564 10500 25620 10668
rect 25564 10434 25620 10444
rect 25228 8932 25284 9772
rect 25228 8866 25284 8876
rect 25340 9604 25396 9614
rect 25340 8930 25396 9548
rect 25452 9042 25508 9884
rect 25452 8990 25454 9042
rect 25506 8990 25508 9042
rect 25452 8978 25508 8990
rect 25564 9154 25620 9166
rect 25564 9102 25566 9154
rect 25618 9102 25620 9154
rect 25340 8878 25342 8930
rect 25394 8878 25396 8930
rect 25340 8596 25396 8878
rect 25340 8530 25396 8540
rect 25452 8820 25508 8830
rect 25228 8372 25284 8382
rect 25228 8148 25284 8316
rect 25228 7586 25284 8092
rect 25228 7534 25230 7586
rect 25282 7534 25284 7586
rect 25228 7522 25284 7534
rect 25340 7588 25396 7598
rect 25340 7494 25396 7532
rect 25340 7252 25396 7262
rect 25340 7158 25396 7196
rect 25228 6020 25284 6030
rect 25228 5926 25284 5964
rect 24892 5234 25060 5236
rect 24892 5182 24894 5234
rect 24946 5182 25060 5234
rect 24892 5180 25060 5182
rect 24892 5170 24948 5180
rect 24780 4510 24782 4562
rect 24834 4510 24836 4562
rect 24780 4498 24836 4510
rect 25228 4452 25284 4462
rect 25452 4452 25508 8764
rect 25228 4450 25508 4452
rect 25228 4398 25230 4450
rect 25282 4398 25508 4450
rect 25228 4396 25508 4398
rect 25228 4386 25284 4396
rect 25564 4228 25620 9102
rect 25676 8932 25732 11900
rect 25900 11284 25956 13806
rect 26124 13636 26180 14590
rect 26124 13580 26292 13636
rect 26124 13300 26180 13310
rect 26124 12962 26180 13244
rect 26236 13074 26292 13580
rect 26236 13022 26238 13074
rect 26290 13022 26292 13074
rect 26236 13010 26292 13022
rect 26124 12910 26126 12962
rect 26178 12910 26180 12962
rect 25900 11218 25956 11228
rect 26012 12290 26068 12302
rect 26012 12238 26014 12290
rect 26066 12238 26068 12290
rect 26012 10722 26068 12238
rect 26124 11732 26180 12910
rect 26236 12850 26292 12862
rect 26236 12798 26238 12850
rect 26290 12798 26292 12850
rect 26236 12178 26292 12798
rect 26236 12126 26238 12178
rect 26290 12126 26292 12178
rect 26236 12114 26292 12126
rect 26124 11666 26180 11676
rect 26124 11396 26180 11406
rect 26124 11302 26180 11340
rect 26012 10670 26014 10722
rect 26066 10670 26068 10722
rect 26012 10658 26068 10670
rect 26236 10610 26292 10622
rect 26236 10558 26238 10610
rect 26290 10558 26292 10610
rect 26236 10388 26292 10558
rect 26236 10322 26292 10332
rect 26348 10052 26404 15092
rect 26572 14418 26628 15036
rect 26572 14366 26574 14418
rect 26626 14366 26628 14418
rect 26572 14354 26628 14366
rect 26908 12964 26964 12974
rect 26908 12870 26964 12908
rect 27020 11508 27076 15260
rect 27132 15148 27188 16828
rect 27468 16882 27524 17164
rect 27580 17108 27636 17390
rect 27692 17444 27748 18510
rect 28140 18450 28196 18732
rect 28140 18398 28142 18450
rect 28194 18398 28196 18450
rect 28140 18340 28196 18398
rect 28140 18274 28196 18284
rect 28252 18004 28308 19180
rect 28588 19124 28644 19516
rect 28476 19068 28644 19124
rect 28364 18564 28420 18574
rect 28364 18470 28420 18508
rect 27692 17378 27748 17388
rect 28140 17948 28308 18004
rect 28140 17778 28196 17948
rect 28140 17726 28142 17778
rect 28194 17726 28196 17778
rect 28140 17444 28196 17726
rect 28140 17378 28196 17388
rect 28252 17780 28308 17790
rect 27916 17108 27972 17118
rect 27580 17106 27972 17108
rect 27580 17054 27918 17106
rect 27970 17054 27972 17106
rect 27580 17052 27972 17054
rect 27468 16830 27470 16882
rect 27522 16830 27524 16882
rect 27468 16660 27524 16830
rect 27356 16604 27524 16660
rect 27580 16772 27636 16782
rect 27356 16548 27412 16604
rect 27580 16548 27636 16716
rect 27356 16482 27412 16492
rect 27468 16492 27636 16548
rect 27468 16100 27524 16492
rect 27468 16006 27524 16044
rect 27580 16324 27636 16334
rect 27580 15986 27636 16268
rect 27580 15934 27582 15986
rect 27634 15934 27636 15986
rect 27356 15540 27412 15550
rect 27356 15426 27412 15484
rect 27356 15374 27358 15426
rect 27410 15374 27412 15426
rect 27356 15362 27412 15374
rect 27580 15148 27636 15934
rect 27692 15764 27748 17052
rect 27916 17042 27972 17052
rect 28140 17108 28196 17118
rect 28252 17108 28308 17724
rect 28140 17106 28308 17108
rect 28140 17054 28142 17106
rect 28194 17054 28308 17106
rect 28140 17052 28308 17054
rect 28140 17042 28196 17052
rect 27804 16884 27860 16894
rect 28364 16884 28420 16894
rect 27804 16790 27860 16828
rect 28252 16882 28420 16884
rect 28252 16830 28366 16882
rect 28418 16830 28420 16882
rect 28252 16828 28420 16830
rect 28252 16324 28308 16828
rect 28364 16818 28420 16828
rect 27916 16268 28308 16324
rect 27916 16210 27972 16268
rect 27916 16158 27918 16210
rect 27970 16158 27972 16210
rect 27916 16146 27972 16158
rect 28140 15876 28196 15886
rect 27692 15708 27860 15764
rect 27692 15316 27748 15326
rect 27692 15222 27748 15260
rect 27132 15092 27524 15148
rect 27580 15092 27748 15148
rect 27356 14644 27412 14654
rect 27132 14420 27188 14430
rect 27132 14326 27188 14364
rect 27356 13748 27412 14588
rect 27468 14532 27524 15092
rect 27468 14438 27524 14476
rect 27580 14980 27636 14990
rect 27356 12962 27412 13692
rect 27580 13634 27636 14924
rect 27692 14868 27748 15092
rect 27804 15092 27860 15708
rect 27804 15026 27860 15036
rect 27692 14812 27860 14868
rect 27692 14420 27748 14430
rect 27692 14084 27748 14364
rect 27692 14018 27748 14028
rect 27580 13582 27582 13634
rect 27634 13582 27636 13634
rect 27580 13570 27636 13582
rect 27692 13748 27748 13758
rect 27804 13748 27860 14812
rect 27916 14418 27972 14430
rect 27916 14366 27918 14418
rect 27970 14366 27972 14418
rect 27916 14196 27972 14366
rect 27916 14130 27972 14140
rect 28028 14306 28084 14318
rect 28028 14254 28030 14306
rect 28082 14254 28084 14306
rect 28028 13972 28084 14254
rect 28028 13906 28084 13916
rect 27692 13746 27860 13748
rect 27692 13694 27694 13746
rect 27746 13694 27860 13746
rect 27692 13692 27860 13694
rect 27692 13412 27748 13692
rect 27356 12910 27358 12962
rect 27410 12910 27412 12962
rect 27356 12898 27412 12910
rect 27468 13356 27748 13412
rect 27132 12740 27188 12750
rect 27132 12178 27188 12684
rect 27132 12126 27134 12178
rect 27186 12126 27188 12178
rect 27132 12114 27188 12126
rect 27356 12178 27412 12190
rect 27356 12126 27358 12178
rect 27410 12126 27412 12178
rect 27356 11844 27412 12126
rect 26908 11452 27076 11508
rect 27132 11788 27412 11844
rect 27132 11506 27188 11788
rect 27132 11454 27134 11506
rect 27186 11454 27188 11506
rect 26684 10612 26740 10622
rect 26684 10518 26740 10556
rect 25676 8866 25732 8876
rect 26124 9996 26404 10052
rect 25788 8260 25844 8270
rect 25788 8166 25844 8204
rect 25788 7700 25844 7710
rect 25676 7644 25788 7700
rect 25676 6244 25732 7644
rect 25788 7634 25844 7644
rect 25900 7476 25956 7486
rect 25900 7474 26068 7476
rect 25900 7422 25902 7474
rect 25954 7422 26068 7474
rect 25900 7420 26068 7422
rect 25900 7410 25956 7420
rect 25676 6188 25956 6244
rect 25788 6020 25844 6030
rect 25116 4172 25564 4228
rect 25116 3666 25172 4172
rect 25564 4134 25620 4172
rect 25676 5964 25788 6020
rect 25676 3780 25732 5964
rect 25788 5954 25844 5964
rect 25900 4452 25956 6188
rect 26012 5684 26068 7420
rect 26012 5122 26068 5628
rect 26012 5070 26014 5122
rect 26066 5070 26068 5122
rect 26012 5058 26068 5070
rect 26124 6578 26180 9996
rect 26236 9828 26292 9838
rect 26684 9828 26740 9838
rect 26236 9826 26740 9828
rect 26236 9774 26238 9826
rect 26290 9774 26686 9826
rect 26738 9774 26740 9826
rect 26236 9772 26740 9774
rect 26236 9762 26292 9772
rect 26684 9156 26740 9772
rect 26684 9090 26740 9100
rect 26460 8932 26516 8942
rect 26236 8596 26292 8606
rect 26236 6690 26292 8540
rect 26348 8148 26404 8158
rect 26348 8054 26404 8092
rect 26348 7588 26404 7598
rect 26460 7588 26516 8876
rect 26908 8484 26964 11452
rect 27132 11442 27188 11454
rect 27244 11394 27300 11406
rect 27244 11342 27246 11394
rect 27298 11342 27300 11394
rect 27020 11284 27076 11294
rect 27020 9828 27076 11228
rect 27244 11284 27300 11342
rect 27244 10052 27300 11228
rect 27244 9986 27300 9996
rect 27356 10050 27412 10062
rect 27356 9998 27358 10050
rect 27410 9998 27412 10050
rect 27356 9940 27412 9998
rect 27356 9874 27412 9884
rect 27020 9734 27076 9772
rect 27132 9044 27188 9054
rect 27132 8950 27188 8988
rect 26908 8418 26964 8428
rect 26348 7586 26516 7588
rect 26348 7534 26350 7586
rect 26402 7534 26516 7586
rect 26348 7532 26516 7534
rect 26348 7522 26404 7532
rect 26236 6638 26238 6690
rect 26290 6638 26292 6690
rect 26236 6626 26292 6638
rect 26124 6526 26126 6578
rect 26178 6526 26180 6578
rect 26124 4900 26180 6526
rect 26124 4834 26180 4844
rect 26236 5906 26292 5918
rect 26236 5854 26238 5906
rect 26290 5854 26292 5906
rect 26236 5572 26292 5854
rect 26460 5796 26516 7532
rect 26796 8034 26852 8046
rect 26796 7982 26798 8034
rect 26850 7982 26852 8034
rect 26460 5730 26516 5740
rect 26572 7028 26628 7038
rect 26572 5684 26628 6972
rect 26684 6804 26740 6814
rect 26796 6804 26852 7982
rect 27020 8036 27076 8046
rect 27244 8036 27300 8046
rect 27076 8034 27300 8036
rect 27076 7982 27246 8034
rect 27298 7982 27300 8034
rect 27076 7980 27300 7982
rect 26740 6748 26964 6804
rect 26684 6738 26740 6748
rect 26684 6468 26740 6478
rect 26684 6374 26740 6412
rect 26908 6468 26964 6748
rect 26908 6402 26964 6412
rect 26796 6132 26852 6142
rect 26796 6038 26852 6076
rect 27020 6020 27076 7980
rect 27244 7970 27300 7980
rect 27244 7474 27300 7486
rect 27244 7422 27246 7474
rect 27298 7422 27300 7474
rect 27244 6804 27300 7422
rect 27356 7028 27412 7038
rect 27468 7028 27524 13356
rect 28140 13300 28196 15820
rect 28252 15428 28308 15438
rect 28252 15334 28308 15372
rect 28476 15148 28532 19068
rect 28812 18564 28868 20412
rect 28924 20412 29372 20468
rect 28924 19572 28980 20412
rect 29372 20374 29428 20412
rect 28924 19506 28980 19516
rect 29036 20018 29092 20030
rect 29036 19966 29038 20018
rect 29090 19966 29092 20018
rect 29036 18676 29092 19966
rect 29260 20020 29316 20030
rect 29260 20018 29428 20020
rect 29260 19966 29262 20018
rect 29314 19966 29428 20018
rect 29260 19964 29428 19966
rect 29260 19954 29316 19964
rect 29148 19906 29204 19918
rect 29148 19854 29150 19906
rect 29202 19854 29204 19906
rect 29148 19236 29204 19854
rect 29260 19236 29316 19246
rect 29148 19234 29316 19236
rect 29148 19182 29262 19234
rect 29314 19182 29316 19234
rect 29148 19180 29316 19182
rect 29260 19170 29316 19180
rect 29036 18610 29092 18620
rect 28924 18564 28980 18574
rect 28812 18508 28924 18564
rect 28700 17442 28756 17454
rect 28700 17390 28702 17442
rect 28754 17390 28756 17442
rect 28588 15874 28644 15886
rect 28588 15822 28590 15874
rect 28642 15822 28644 15874
rect 28588 15764 28644 15822
rect 28588 15698 28644 15708
rect 28252 15092 28532 15148
rect 28588 15428 28644 15438
rect 28588 15148 28644 15372
rect 28700 15316 28756 17390
rect 28924 16324 28980 18508
rect 29036 18450 29092 18462
rect 29036 18398 29038 18450
rect 29090 18398 29092 18450
rect 29036 18228 29092 18398
rect 29036 18162 29092 18172
rect 29372 17668 29428 19964
rect 29484 19684 29540 23660
rect 30268 23716 30324 23774
rect 30268 23650 30324 23660
rect 30604 23716 30660 23726
rect 30604 23622 30660 23660
rect 30716 23714 30772 24108
rect 30716 23662 30718 23714
rect 30770 23662 30772 23714
rect 29596 23154 29652 23166
rect 29596 23102 29598 23154
rect 29650 23102 29652 23154
rect 29596 20916 29652 23102
rect 29932 23154 29988 23166
rect 29932 23102 29934 23154
rect 29986 23102 29988 23154
rect 29932 22372 29988 23102
rect 30380 23154 30436 23166
rect 30380 23102 30382 23154
rect 30434 23102 30436 23154
rect 30380 23044 30436 23102
rect 30044 22930 30100 22942
rect 30044 22878 30046 22930
rect 30098 22878 30100 22930
rect 30044 22482 30100 22878
rect 30044 22430 30046 22482
rect 30098 22430 30100 22482
rect 30044 22418 30100 22430
rect 30268 22932 30324 22942
rect 29932 22306 29988 22316
rect 30268 22370 30324 22876
rect 30268 22318 30270 22370
rect 30322 22318 30324 22370
rect 30268 22306 30324 22318
rect 30044 22260 30100 22270
rect 29708 22148 29764 22158
rect 29708 21586 29764 22092
rect 29708 21534 29710 21586
rect 29762 21534 29764 21586
rect 29708 21522 29764 21534
rect 30044 21474 30100 22204
rect 30044 21422 30046 21474
rect 30098 21422 30100 21474
rect 30044 21410 30100 21422
rect 30156 21586 30212 21598
rect 30156 21534 30158 21586
rect 30210 21534 30212 21586
rect 30156 21028 30212 21534
rect 30156 20962 30212 20972
rect 30268 21476 30324 21486
rect 30268 21026 30324 21420
rect 30268 20974 30270 21026
rect 30322 20974 30324 21026
rect 30268 20962 30324 20974
rect 29596 20850 29652 20860
rect 30156 20690 30212 20702
rect 30156 20638 30158 20690
rect 30210 20638 30212 20690
rect 29932 20580 29988 20590
rect 29932 20486 29988 20524
rect 29708 20018 29764 20030
rect 29708 19966 29710 20018
rect 29762 19966 29764 20018
rect 29708 19908 29764 19966
rect 30156 20020 30212 20638
rect 30268 20578 30324 20590
rect 30268 20526 30270 20578
rect 30322 20526 30324 20578
rect 30268 20244 30324 20526
rect 30380 20580 30436 22988
rect 30716 22036 30772 23662
rect 30940 23938 30996 23950
rect 30940 23886 30942 23938
rect 30994 23886 30996 23938
rect 30940 23154 30996 23886
rect 30940 23102 30942 23154
rect 30994 23102 30996 23154
rect 30940 22260 30996 23102
rect 31052 22932 31108 24558
rect 31164 23940 31220 24668
rect 31276 24630 31332 24668
rect 31164 23874 31220 23884
rect 31724 24610 31780 24622
rect 31724 24558 31726 24610
rect 31778 24558 31780 24610
rect 31724 23938 31780 24558
rect 31724 23886 31726 23938
rect 31778 23886 31780 23938
rect 31724 23604 31780 23886
rect 31836 23826 31892 25116
rect 31836 23774 31838 23826
rect 31890 23774 31892 23826
rect 31836 23762 31892 23774
rect 31948 25060 32004 25070
rect 31724 23538 31780 23548
rect 31836 23268 31892 23278
rect 31052 22866 31108 22876
rect 31388 23154 31444 23166
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 31388 22708 31444 23102
rect 31500 23156 31556 23166
rect 31500 23062 31556 23100
rect 31612 23156 31668 23166
rect 31836 23156 31892 23212
rect 31612 23154 31892 23156
rect 31612 23102 31614 23154
rect 31666 23102 31892 23154
rect 31612 23100 31892 23102
rect 31612 23090 31668 23100
rect 31388 22642 31444 22652
rect 31276 22596 31332 22606
rect 31276 22502 31332 22540
rect 30940 22194 30996 22204
rect 31052 22482 31108 22494
rect 31052 22430 31054 22482
rect 31106 22430 31108 22482
rect 30716 21970 30772 21980
rect 30828 21588 30884 21598
rect 30828 21494 30884 21532
rect 31052 21586 31108 22430
rect 31388 22370 31444 22382
rect 31388 22318 31390 22370
rect 31442 22318 31444 22370
rect 31388 21700 31444 22318
rect 31444 21644 31668 21700
rect 31388 21634 31444 21644
rect 31052 21534 31054 21586
rect 31106 21534 31108 21586
rect 31052 21476 31108 21534
rect 31052 21410 31108 21420
rect 31276 21364 31332 21374
rect 31276 21270 31332 21308
rect 30380 20514 30436 20524
rect 30828 21028 30884 21038
rect 30268 20178 30324 20188
rect 30492 20356 30548 20366
rect 30380 20020 30436 20030
rect 30156 20018 30436 20020
rect 30156 19966 30382 20018
rect 30434 19966 30436 20018
rect 30156 19964 30436 19966
rect 30044 19908 30100 19918
rect 29708 19906 30100 19908
rect 29708 19854 30046 19906
rect 30098 19854 30100 19906
rect 29708 19852 30100 19854
rect 30044 19796 30100 19852
rect 30156 19796 30212 19806
rect 30044 19740 30156 19796
rect 30156 19730 30212 19740
rect 29484 19628 30100 19684
rect 29484 19236 29540 19246
rect 29484 19142 29540 19180
rect 29596 18676 29652 18686
rect 29596 18582 29652 18620
rect 29820 18226 29876 18238
rect 29820 18174 29822 18226
rect 29874 18174 29876 18226
rect 29260 17612 29428 17668
rect 29596 17666 29652 17678
rect 29596 17614 29598 17666
rect 29650 17614 29652 17666
rect 28924 16258 28980 16268
rect 29036 17444 29092 17454
rect 28812 15988 28868 15998
rect 28812 15538 28868 15932
rect 28812 15486 28814 15538
rect 28866 15486 28868 15538
rect 28812 15474 28868 15486
rect 28700 15250 28756 15260
rect 29036 15148 29092 17388
rect 29148 16996 29204 17006
rect 29148 16882 29204 16940
rect 29148 16830 29150 16882
rect 29202 16830 29204 16882
rect 29148 16818 29204 16830
rect 29148 16548 29204 16558
rect 29148 15426 29204 16492
rect 29260 16436 29316 17612
rect 29372 17442 29428 17454
rect 29372 17390 29374 17442
rect 29426 17390 29428 17442
rect 29372 17108 29428 17390
rect 29596 17220 29652 17614
rect 29596 17154 29652 17164
rect 29372 17042 29428 17052
rect 29484 16772 29540 16782
rect 29820 16772 29876 18174
rect 29484 16770 29876 16772
rect 29484 16718 29486 16770
rect 29538 16718 29876 16770
rect 29484 16716 29876 16718
rect 29932 17108 29988 17118
rect 29484 16706 29540 16716
rect 29372 16492 29652 16548
rect 29372 16436 29428 16492
rect 29260 16380 29428 16436
rect 29148 15374 29150 15426
rect 29202 15374 29204 15426
rect 29148 15362 29204 15374
rect 29484 16324 29540 16334
rect 29372 15316 29428 15326
rect 29260 15314 29428 15316
rect 29260 15262 29374 15314
rect 29426 15262 29428 15314
rect 29260 15260 29428 15262
rect 29260 15148 29316 15260
rect 29372 15250 29428 15260
rect 28588 15092 28756 15148
rect 28252 14532 28308 15092
rect 28588 14980 28644 14990
rect 28588 14642 28644 14924
rect 28588 14590 28590 14642
rect 28642 14590 28644 14642
rect 28588 14578 28644 14590
rect 28252 14466 28308 14476
rect 28476 14532 28532 14542
rect 28252 14308 28308 14318
rect 28252 14306 28420 14308
rect 28252 14254 28254 14306
rect 28306 14254 28420 14306
rect 28252 14252 28420 14254
rect 28252 14242 28308 14252
rect 28364 13746 28420 14252
rect 28364 13694 28366 13746
rect 28418 13694 28420 13746
rect 28364 13682 28420 13694
rect 28476 13524 28532 14476
rect 27580 13244 28196 13300
rect 28252 13300 28308 13310
rect 27580 11508 27636 13244
rect 28252 13076 28308 13244
rect 28028 12964 28084 12974
rect 28252 12964 28308 13020
rect 28028 12962 28308 12964
rect 28028 12910 28030 12962
rect 28082 12910 28308 12962
rect 28028 12908 28308 12910
rect 28364 12964 28420 12974
rect 28476 12964 28532 13468
rect 28364 12962 28532 12964
rect 28364 12910 28366 12962
rect 28418 12910 28532 12962
rect 28364 12908 28532 12910
rect 28588 12964 28644 12974
rect 28700 12964 28756 15092
rect 29036 15092 29316 15148
rect 28588 12962 28756 12964
rect 28588 12910 28590 12962
rect 28642 12910 28756 12962
rect 28588 12908 28756 12910
rect 28924 14196 28980 14206
rect 28924 13746 28980 14140
rect 28924 13694 28926 13746
rect 28978 13694 28980 13746
rect 28028 12898 28084 12908
rect 28364 12898 28420 12908
rect 28028 12740 28084 12750
rect 27580 11442 27636 11452
rect 27804 12516 27860 12526
rect 27804 11394 27860 12460
rect 27804 11342 27806 11394
rect 27858 11342 27860 11394
rect 27804 11330 27860 11342
rect 28028 11172 28084 12684
rect 27692 11116 28084 11172
rect 28140 12738 28196 12750
rect 28140 12686 28142 12738
rect 28194 12686 28196 12738
rect 27580 10836 27636 10846
rect 27580 10742 27636 10780
rect 27692 9604 27748 11116
rect 28140 10724 28196 12686
rect 28252 12738 28308 12750
rect 28252 12686 28254 12738
rect 28306 12686 28308 12738
rect 28252 12068 28308 12686
rect 28252 12002 28308 12012
rect 28364 11956 28420 11966
rect 28364 11862 28420 11900
rect 28588 11732 28644 12908
rect 28588 11666 28644 11676
rect 28700 11620 28756 11630
rect 28028 10668 28196 10724
rect 28252 11394 28308 11406
rect 28252 11342 28254 11394
rect 28306 11342 28308 11394
rect 27916 10052 27972 10062
rect 28028 10052 28084 10668
rect 28140 10500 28196 10510
rect 28140 10406 28196 10444
rect 28252 10052 28308 11342
rect 28364 11282 28420 11294
rect 28364 11230 28366 11282
rect 28418 11230 28420 11282
rect 28364 10836 28420 11230
rect 28700 11284 28756 11564
rect 28700 11218 28756 11228
rect 28364 10770 28420 10780
rect 28588 10722 28644 10734
rect 28588 10670 28590 10722
rect 28642 10670 28644 10722
rect 28364 10052 28420 10062
rect 28028 9996 28196 10052
rect 28252 10050 28420 10052
rect 28252 9998 28366 10050
rect 28418 9998 28420 10050
rect 28252 9996 28420 9998
rect 27916 9940 27972 9996
rect 27916 9884 28084 9940
rect 27804 9826 27860 9838
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9716 27860 9774
rect 28028 9826 28084 9884
rect 28028 9774 28030 9826
rect 28082 9774 28084 9826
rect 28028 9762 28084 9774
rect 27804 9660 27972 9716
rect 27692 9548 27860 9604
rect 27692 9268 27748 9278
rect 27412 6972 27524 7028
rect 27580 9212 27692 9268
rect 27356 6962 27412 6972
rect 27580 6804 27636 9212
rect 27692 9174 27748 9212
rect 27692 8258 27748 8270
rect 27692 8206 27694 8258
rect 27746 8206 27748 8258
rect 27692 7812 27748 8206
rect 27692 7140 27748 7756
rect 27804 7362 27860 9548
rect 27916 7700 27972 9660
rect 28140 9604 28196 9996
rect 28364 9986 28420 9996
rect 28252 9828 28308 9838
rect 28252 9734 28308 9772
rect 28140 9548 28308 9604
rect 28028 9156 28084 9166
rect 28028 9062 28084 9100
rect 28028 8260 28084 8270
rect 28028 7924 28084 8204
rect 28028 7858 28084 7868
rect 28140 8146 28196 8158
rect 28140 8094 28142 8146
rect 28194 8094 28196 8146
rect 27916 7634 27972 7644
rect 28140 7700 28196 8094
rect 28028 7588 28084 7598
rect 27804 7310 27806 7362
rect 27858 7310 27860 7362
rect 27804 7298 27860 7310
rect 27916 7476 27972 7486
rect 27916 7140 27972 7420
rect 27692 7084 27860 7140
rect 27020 5954 27076 5964
rect 27132 6748 27244 6804
rect 27132 5796 27188 6748
rect 27244 6738 27300 6748
rect 27356 6748 27636 6804
rect 27692 6916 27748 6926
rect 27244 6468 27300 6478
rect 27244 6374 27300 6412
rect 27356 6018 27412 6748
rect 27356 5966 27358 6018
rect 27410 5966 27412 6018
rect 27356 5908 27412 5966
rect 27356 5842 27412 5852
rect 27468 6468 27524 6478
rect 26908 5740 27188 5796
rect 27244 5794 27300 5806
rect 27244 5742 27246 5794
rect 27298 5742 27300 5794
rect 26572 5628 26852 5684
rect 26236 4564 26292 5516
rect 26348 5348 26404 5358
rect 26348 5010 26404 5292
rect 26572 5236 26628 5246
rect 26572 5142 26628 5180
rect 26348 4958 26350 5010
rect 26402 4958 26404 5010
rect 26348 4900 26404 4958
rect 26572 5012 26628 5022
rect 26348 4834 26404 4844
rect 26460 4898 26516 4910
rect 26460 4846 26462 4898
rect 26514 4846 26516 4898
rect 26236 4498 26292 4508
rect 25900 4396 26180 4452
rect 25788 4340 25844 4350
rect 25788 4338 25956 4340
rect 25788 4286 25790 4338
rect 25842 4286 25956 4338
rect 25788 4284 25956 4286
rect 25788 4274 25844 4284
rect 25788 3780 25844 3790
rect 25676 3778 25844 3780
rect 25676 3726 25790 3778
rect 25842 3726 25844 3778
rect 25676 3724 25844 3726
rect 25788 3714 25844 3724
rect 25116 3614 25118 3666
rect 25170 3614 25172 3666
rect 25116 3602 25172 3614
rect 25900 3556 25956 4284
rect 26124 3778 26180 4396
rect 26124 3726 26126 3778
rect 26178 3726 26180 3778
rect 26124 3714 26180 3726
rect 26460 4338 26516 4846
rect 26460 4286 26462 4338
rect 26514 4286 26516 4338
rect 26124 3556 26180 3566
rect 26460 3556 26516 4286
rect 25900 3554 26516 3556
rect 25900 3502 26126 3554
rect 26178 3502 26516 3554
rect 25900 3500 26516 3502
rect 26572 3556 26628 4956
rect 26684 4898 26740 4910
rect 26684 4846 26686 4898
rect 26738 4846 26740 4898
rect 26684 4340 26740 4846
rect 26684 4274 26740 4284
rect 26796 4226 26852 5628
rect 26796 4174 26798 4226
rect 26850 4174 26852 4226
rect 26796 4162 26852 4174
rect 26684 3556 26740 3566
rect 26572 3554 26740 3556
rect 26572 3502 26686 3554
rect 26738 3502 26740 3554
rect 26572 3500 26740 3502
rect 26124 3490 26180 3500
rect 26460 3442 26516 3500
rect 26684 3490 26740 3500
rect 26460 3390 26462 3442
rect 26514 3390 26516 3442
rect 26460 3378 26516 3390
rect 24668 2258 24724 2268
rect 18844 1586 18900 1596
rect 26908 1652 26964 5740
rect 27132 5236 27188 5246
rect 27244 5236 27300 5742
rect 27132 5234 27300 5236
rect 27132 5182 27134 5234
rect 27186 5182 27300 5234
rect 27132 5180 27300 5182
rect 27356 5236 27412 5246
rect 27132 5170 27188 5180
rect 27356 5142 27412 5180
rect 27356 4900 27412 4910
rect 27244 4564 27300 4574
rect 27244 4470 27300 4508
rect 27356 3668 27412 4844
rect 27468 4564 27524 6412
rect 27692 6132 27748 6860
rect 27804 6802 27860 7084
rect 27916 7074 27972 7084
rect 27804 6750 27806 6802
rect 27858 6750 27860 6802
rect 27804 6580 27860 6750
rect 27804 6514 27860 6524
rect 27804 6132 27860 6142
rect 27692 6130 27860 6132
rect 27692 6078 27806 6130
rect 27858 6078 27860 6130
rect 27692 6076 27860 6078
rect 27804 6066 27860 6076
rect 27580 6020 27636 6030
rect 27580 5926 27636 5964
rect 27804 5908 27860 5918
rect 27692 5684 27748 5694
rect 27692 5346 27748 5628
rect 27692 5294 27694 5346
rect 27746 5294 27748 5346
rect 27692 5282 27748 5294
rect 27468 4498 27524 4508
rect 27804 4338 27860 5852
rect 28028 4564 28084 7532
rect 28140 7476 28196 7644
rect 28140 7410 28196 7420
rect 28140 7252 28196 7262
rect 28140 5906 28196 7196
rect 28252 6690 28308 9548
rect 28588 9042 28644 10670
rect 28812 10610 28868 10622
rect 28812 10558 28814 10610
rect 28866 10558 28868 10610
rect 28588 8990 28590 9042
rect 28642 8990 28644 9042
rect 28588 8978 28644 8990
rect 28700 10498 28756 10510
rect 28700 10446 28702 10498
rect 28754 10446 28756 10498
rect 28700 9828 28756 10446
rect 28700 8428 28756 9772
rect 28812 9268 28868 10558
rect 28924 10500 28980 13694
rect 28924 10434 28980 10444
rect 28812 9202 28868 9212
rect 29036 8596 29092 15092
rect 29148 14308 29204 14318
rect 29148 14214 29204 14252
rect 29372 14084 29428 14094
rect 29260 13522 29316 13534
rect 29260 13470 29262 13522
rect 29314 13470 29316 13522
rect 29260 12962 29316 13470
rect 29260 12910 29262 12962
rect 29314 12910 29316 12962
rect 29260 12898 29316 12910
rect 29372 11956 29428 14028
rect 29484 12178 29540 16268
rect 29484 12126 29486 12178
rect 29538 12126 29540 12178
rect 29484 12114 29540 12126
rect 29372 11900 29540 11956
rect 29484 11394 29540 11900
rect 29484 11342 29486 11394
rect 29538 11342 29540 11394
rect 29484 11330 29540 11342
rect 29260 11282 29316 11294
rect 29260 11230 29262 11282
rect 29314 11230 29316 11282
rect 29148 10948 29204 10958
rect 29260 10948 29316 11230
rect 29204 10892 29316 10948
rect 29148 10882 29204 10892
rect 28252 6638 28254 6690
rect 28306 6638 28308 6690
rect 28252 6626 28308 6638
rect 28364 8372 28420 8382
rect 28140 5854 28142 5906
rect 28194 5854 28196 5906
rect 28140 5122 28196 5854
rect 28252 5682 28308 5694
rect 28252 5630 28254 5682
rect 28306 5630 28308 5682
rect 28252 5572 28308 5630
rect 28252 5506 28308 5516
rect 28364 5236 28420 8316
rect 28476 8370 28532 8382
rect 28476 8318 28478 8370
rect 28530 8318 28532 8370
rect 28476 7252 28532 8318
rect 28588 8372 28756 8428
rect 28924 8540 29092 8596
rect 29148 9156 29204 9166
rect 28588 7588 28644 8372
rect 28588 7522 28644 7532
rect 28476 7186 28532 7196
rect 28588 6580 28644 6590
rect 28812 6580 28868 6590
rect 28588 6578 28756 6580
rect 28588 6526 28590 6578
rect 28642 6526 28756 6578
rect 28588 6524 28756 6526
rect 28588 6514 28644 6524
rect 28476 6466 28532 6478
rect 28476 6414 28478 6466
rect 28530 6414 28532 6466
rect 28476 5796 28532 6414
rect 28476 5460 28532 5740
rect 28476 5404 28644 5460
rect 28476 5236 28532 5246
rect 28364 5234 28532 5236
rect 28364 5182 28478 5234
rect 28530 5182 28532 5234
rect 28364 5180 28532 5182
rect 28476 5170 28532 5180
rect 28140 5070 28142 5122
rect 28194 5070 28196 5122
rect 28140 5058 28196 5070
rect 28588 5012 28644 5404
rect 28476 4956 28644 5012
rect 28364 4564 28420 4574
rect 28028 4562 28420 4564
rect 28028 4510 28366 4562
rect 28418 4510 28420 4562
rect 28028 4508 28420 4510
rect 28364 4498 28420 4508
rect 27804 4286 27806 4338
rect 27858 4286 27860 4338
rect 27804 4274 27860 4286
rect 27356 3574 27412 3612
rect 27804 3556 27860 3566
rect 27804 3462 27860 3500
rect 28476 3556 28532 4956
rect 28588 4788 28644 4798
rect 28588 4338 28644 4732
rect 28588 4286 28590 4338
rect 28642 4286 28644 4338
rect 28588 4274 28644 4286
rect 28700 4228 28756 6524
rect 28812 5906 28868 6524
rect 28812 5854 28814 5906
rect 28866 5854 28868 5906
rect 28812 5842 28868 5854
rect 28924 4788 28980 8540
rect 29036 8148 29092 8158
rect 29036 7362 29092 8092
rect 29148 7476 29204 9100
rect 29260 9044 29316 10892
rect 29372 11282 29428 11294
rect 29372 11230 29374 11282
rect 29426 11230 29428 11282
rect 29372 11172 29428 11230
rect 29596 11172 29652 16492
rect 29932 16436 29988 17052
rect 29820 16380 29988 16436
rect 29820 16098 29876 16380
rect 30044 16324 30100 19628
rect 30268 19236 30324 19964
rect 30380 19954 30436 19964
rect 30380 19460 30436 19470
rect 30380 19366 30436 19404
rect 30156 19180 30324 19236
rect 30492 19234 30548 20300
rect 30492 19182 30494 19234
rect 30546 19182 30548 19234
rect 30156 16996 30212 19180
rect 30492 19170 30548 19182
rect 30604 19684 30660 19694
rect 30268 19012 30324 19022
rect 30268 18450 30324 18956
rect 30268 18398 30270 18450
rect 30322 18398 30324 18450
rect 30268 18386 30324 18398
rect 30380 18450 30436 18462
rect 30380 18398 30382 18450
rect 30434 18398 30436 18450
rect 30380 17892 30436 18398
rect 30380 17826 30436 17836
rect 30492 18452 30548 18462
rect 30492 17890 30548 18396
rect 30492 17838 30494 17890
rect 30546 17838 30548 17890
rect 30156 16930 30212 16940
rect 30268 17220 30324 17230
rect 29820 16046 29822 16098
rect 29874 16046 29876 16098
rect 29820 14644 29876 16046
rect 29932 16268 30100 16324
rect 29932 15764 29988 16268
rect 29932 15148 29988 15708
rect 30044 15986 30100 15998
rect 30044 15934 30046 15986
rect 30098 15934 30100 15986
rect 30044 15426 30100 15934
rect 30044 15374 30046 15426
rect 30098 15374 30100 15426
rect 30044 15362 30100 15374
rect 30156 15428 30212 15438
rect 30156 15334 30212 15372
rect 29932 15092 30100 15148
rect 29820 14578 29876 14588
rect 29708 14530 29764 14542
rect 29708 14478 29710 14530
rect 29762 14478 29764 14530
rect 29708 14420 29764 14478
rect 29708 14354 29764 14364
rect 29820 12180 29876 12190
rect 29820 12086 29876 12124
rect 29708 12068 29764 12078
rect 29708 11974 29764 12012
rect 29372 11116 29652 11172
rect 29820 11732 29876 11742
rect 29372 10612 29428 11116
rect 29372 10546 29428 10556
rect 29820 10610 29876 11676
rect 29820 10558 29822 10610
rect 29874 10558 29876 10610
rect 29820 10276 29876 10558
rect 29820 10210 29876 10220
rect 29932 11170 29988 11182
rect 29932 11118 29934 11170
rect 29986 11118 29988 11170
rect 29596 9826 29652 9838
rect 29596 9774 29598 9826
rect 29650 9774 29652 9826
rect 29596 9266 29652 9774
rect 29932 9826 29988 11118
rect 29932 9774 29934 9826
rect 29986 9774 29988 9826
rect 29932 9762 29988 9774
rect 29596 9214 29598 9266
rect 29650 9214 29652 9266
rect 29596 9202 29652 9214
rect 29820 9044 29876 9054
rect 29260 9042 29876 9044
rect 29260 8990 29822 9042
rect 29874 8990 29876 9042
rect 29260 8988 29876 8990
rect 29372 8260 29428 8270
rect 29372 8166 29428 8204
rect 29148 7382 29204 7420
rect 29036 7310 29038 7362
rect 29090 7310 29092 7362
rect 29036 6916 29092 7310
rect 29036 6860 29540 6916
rect 29484 6802 29540 6860
rect 29484 6750 29486 6802
rect 29538 6750 29540 6802
rect 29484 6738 29540 6750
rect 29372 6690 29428 6702
rect 29372 6638 29374 6690
rect 29426 6638 29428 6690
rect 29148 5908 29204 5918
rect 28924 4722 28980 4732
rect 29036 5124 29092 5134
rect 28700 4162 28756 4172
rect 28588 3778 28644 3790
rect 28588 3726 28590 3778
rect 28642 3726 28644 3778
rect 28588 3666 28644 3726
rect 28588 3614 28590 3666
rect 28642 3614 28644 3666
rect 28588 3602 28644 3614
rect 29036 3666 29092 5068
rect 29148 5122 29204 5852
rect 29148 5070 29150 5122
rect 29202 5070 29204 5122
rect 29148 5058 29204 5070
rect 29260 5012 29316 5022
rect 29148 4564 29204 4574
rect 29260 4564 29316 4956
rect 29148 4562 29316 4564
rect 29148 4510 29150 4562
rect 29202 4510 29316 4562
rect 29148 4508 29316 4510
rect 29148 4340 29204 4508
rect 29372 4340 29428 6638
rect 29484 4340 29540 4350
rect 29372 4338 29540 4340
rect 29372 4286 29486 4338
rect 29538 4286 29540 4338
rect 29372 4284 29540 4286
rect 29148 4274 29204 4284
rect 29484 4228 29540 4284
rect 29484 4162 29540 4172
rect 29484 3780 29540 3790
rect 29596 3780 29652 8988
rect 29820 8978 29876 8988
rect 29708 8484 29764 8494
rect 29708 6020 29764 8428
rect 30044 8372 30100 15092
rect 30156 14980 30212 14990
rect 30156 14530 30212 14924
rect 30156 14478 30158 14530
rect 30210 14478 30212 14530
rect 30156 14466 30212 14478
rect 30268 13970 30324 17164
rect 30492 17108 30548 17838
rect 30604 18450 30660 19628
rect 30604 18398 30606 18450
rect 30658 18398 30660 18450
rect 30604 17778 30660 18398
rect 30604 17726 30606 17778
rect 30658 17726 30660 17778
rect 30604 17714 30660 17726
rect 30828 19346 30884 20972
rect 31164 20802 31220 20814
rect 31164 20750 31166 20802
rect 31218 20750 31220 20802
rect 31164 20692 31220 20750
rect 31164 20244 31220 20636
rect 31388 20802 31444 20814
rect 31388 20750 31390 20802
rect 31442 20750 31444 20802
rect 31388 20580 31444 20750
rect 31612 20690 31668 21644
rect 31724 21140 31780 21150
rect 31724 20914 31780 21084
rect 31724 20862 31726 20914
rect 31778 20862 31780 20914
rect 31724 20850 31780 20862
rect 31612 20638 31614 20690
rect 31666 20638 31668 20690
rect 31612 20626 31668 20638
rect 31388 20468 31444 20524
rect 31164 20178 31220 20188
rect 31276 20412 31444 20468
rect 31836 20578 31892 23100
rect 31948 21028 32004 25004
rect 32060 24724 32116 24734
rect 32060 24630 32116 24668
rect 32620 24612 32676 24622
rect 32508 23268 32564 23278
rect 32508 23174 32564 23212
rect 32172 23044 32228 23054
rect 32172 22950 32228 22988
rect 32508 22708 32564 22718
rect 32396 21698 32452 21710
rect 32396 21646 32398 21698
rect 32450 21646 32452 21698
rect 32284 21586 32340 21598
rect 32284 21534 32286 21586
rect 32338 21534 32340 21586
rect 32284 21140 32340 21534
rect 32284 21074 32340 21084
rect 31948 20972 32116 21028
rect 31836 20526 31838 20578
rect 31890 20526 31892 20578
rect 31836 20468 31892 20526
rect 30828 19294 30830 19346
rect 30882 19294 30884 19346
rect 30716 17668 30772 17678
rect 30716 17574 30772 17612
rect 30828 17444 30884 19294
rect 30940 19908 30996 19918
rect 30940 18116 30996 19852
rect 30940 18050 30996 18060
rect 31052 18338 31108 18350
rect 31052 18286 31054 18338
rect 31106 18286 31108 18338
rect 31052 17892 31108 18286
rect 31052 17826 31108 17836
rect 30492 17042 30548 17052
rect 30716 17388 30884 17444
rect 30940 17556 30996 17566
rect 30380 15540 30436 15550
rect 30380 15314 30436 15484
rect 30380 15262 30382 15314
rect 30434 15262 30436 15314
rect 30380 15250 30436 15262
rect 30268 13918 30270 13970
rect 30322 13918 30324 13970
rect 30268 13906 30324 13918
rect 30268 13076 30324 13086
rect 30044 8306 30100 8316
rect 30156 13020 30268 13076
rect 29932 8260 29988 8270
rect 29932 8166 29988 8204
rect 30156 7812 30212 13020
rect 30268 13010 30324 13020
rect 30380 12962 30436 12974
rect 30380 12910 30382 12962
rect 30434 12910 30436 12962
rect 30380 12290 30436 12910
rect 30716 12964 30772 17388
rect 30828 16996 30884 17006
rect 30828 16098 30884 16940
rect 30828 16046 30830 16098
rect 30882 16046 30884 16098
rect 30828 13858 30884 16046
rect 30940 15986 30996 17500
rect 30940 15934 30942 15986
rect 30994 15934 30996 15986
rect 30940 15922 30996 15934
rect 31052 17108 31108 17118
rect 31052 15148 31108 17052
rect 31276 16100 31332 20412
rect 31836 20402 31892 20412
rect 31836 20132 31892 20142
rect 31500 19236 31556 19246
rect 31500 19142 31556 19180
rect 31724 17668 31780 17678
rect 31500 17442 31556 17454
rect 31500 17390 31502 17442
rect 31554 17390 31556 17442
rect 31388 16882 31444 16894
rect 31388 16830 31390 16882
rect 31442 16830 31444 16882
rect 31388 16322 31444 16830
rect 31500 16884 31556 17390
rect 31500 16818 31556 16828
rect 31388 16270 31390 16322
rect 31442 16270 31444 16322
rect 31388 16258 31444 16270
rect 31276 16044 31444 16100
rect 31164 15764 31220 15774
rect 31164 15314 31220 15708
rect 31164 15262 31166 15314
rect 31218 15262 31220 15314
rect 31164 15250 31220 15262
rect 31388 15148 31444 16044
rect 31612 15426 31668 15438
rect 31612 15374 31614 15426
rect 31666 15374 31668 15426
rect 31052 15092 31220 15148
rect 30828 13806 30830 13858
rect 30882 13806 30884 13858
rect 30828 13794 30884 13806
rect 31052 13748 31108 13758
rect 31052 13654 31108 13692
rect 30716 12898 30772 12908
rect 30828 13636 30884 13646
rect 30380 12238 30382 12290
rect 30434 12238 30436 12290
rect 30380 12226 30436 12238
rect 30716 12178 30772 12190
rect 30716 12126 30718 12178
rect 30770 12126 30772 12178
rect 30716 11508 30772 12126
rect 30828 11618 30884 13580
rect 30828 11566 30830 11618
rect 30882 11566 30884 11618
rect 30828 11554 30884 11566
rect 31052 13524 31108 13534
rect 30380 11452 30772 11508
rect 30268 10612 30324 10622
rect 30268 10518 30324 10556
rect 30380 8036 30436 11452
rect 30828 11396 30884 11406
rect 31052 11396 31108 13468
rect 30828 11394 31108 11396
rect 30828 11342 30830 11394
rect 30882 11342 31108 11394
rect 30828 11340 31108 11342
rect 30828 11330 30884 11340
rect 30492 11284 30548 11294
rect 30716 11284 30772 11294
rect 30492 11190 30548 11228
rect 30604 11228 30716 11284
rect 30604 8372 30660 11228
rect 30716 11218 30772 11228
rect 31052 10724 31108 10734
rect 30716 10500 30772 10510
rect 30828 10500 30884 10510
rect 30716 10498 30828 10500
rect 30716 10446 30718 10498
rect 30770 10446 30828 10498
rect 30716 10444 30828 10446
rect 30716 10434 30772 10444
rect 30604 8306 30660 8316
rect 30604 8148 30660 8158
rect 30380 7942 30436 7980
rect 30492 8092 30604 8148
rect 29932 7756 30212 7812
rect 29932 6692 29988 7756
rect 30156 7588 30212 7598
rect 29932 6690 30100 6692
rect 29932 6638 29934 6690
rect 29986 6638 30100 6690
rect 29932 6636 30100 6638
rect 29932 6626 29988 6636
rect 29708 5124 29764 5964
rect 29932 5906 29988 5918
rect 29932 5854 29934 5906
rect 29986 5854 29988 5906
rect 29932 5348 29988 5854
rect 30044 5794 30100 6636
rect 30156 6018 30212 7532
rect 30380 7476 30436 7486
rect 30380 7382 30436 7420
rect 30156 5966 30158 6018
rect 30210 5966 30212 6018
rect 30156 5954 30212 5966
rect 30044 5742 30046 5794
rect 30098 5742 30100 5794
rect 30044 5730 30100 5742
rect 29932 5282 29988 5292
rect 29708 4228 29764 5068
rect 30044 5012 30100 5022
rect 30044 4918 30100 4956
rect 30492 4340 30548 8092
rect 30604 8054 30660 8092
rect 30828 8146 30884 10444
rect 30940 9044 30996 9054
rect 30940 8370 30996 8988
rect 30940 8318 30942 8370
rect 30994 8318 30996 8370
rect 30940 8306 30996 8318
rect 30828 8094 30830 8146
rect 30882 8094 30884 8146
rect 30828 8082 30884 8094
rect 30940 8036 30996 8046
rect 30716 7700 30772 7710
rect 30716 7476 30772 7644
rect 30716 7362 30772 7420
rect 30828 7476 30884 7486
rect 30940 7476 30996 7980
rect 31052 7812 31108 10668
rect 31164 9828 31220 15092
rect 31276 15090 31332 15102
rect 31388 15092 31556 15148
rect 31276 15038 31278 15090
rect 31330 15038 31332 15090
rect 31276 14756 31332 15038
rect 31276 14690 31332 14700
rect 31388 14644 31444 14654
rect 31276 14532 31332 14542
rect 31276 14438 31332 14476
rect 31388 13188 31444 14588
rect 31276 13132 31444 13188
rect 31276 11508 31332 13132
rect 31388 12964 31444 12974
rect 31388 12870 31444 12908
rect 31388 12740 31444 12750
rect 31388 12646 31444 12684
rect 31388 12292 31444 12302
rect 31388 12066 31444 12236
rect 31388 12014 31390 12066
rect 31442 12014 31444 12066
rect 31388 12002 31444 12014
rect 31388 11508 31444 11518
rect 31276 11506 31444 11508
rect 31276 11454 31390 11506
rect 31442 11454 31444 11506
rect 31276 11452 31444 11454
rect 31388 11442 31444 11452
rect 31388 10948 31444 10958
rect 31388 10610 31444 10892
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 31388 10546 31444 10558
rect 31500 10388 31556 15092
rect 31612 14196 31668 15374
rect 31612 14130 31668 14140
rect 31724 14420 31780 17612
rect 31836 17556 31892 20076
rect 32060 19460 32116 20972
rect 32396 20244 32452 21646
rect 32284 20188 32452 20244
rect 32172 19908 32228 19918
rect 32284 19908 32340 20188
rect 32396 20020 32452 20030
rect 32396 19926 32452 19964
rect 32228 19852 32340 19908
rect 32172 19842 32228 19852
rect 32060 19394 32116 19404
rect 31948 19346 32004 19358
rect 31948 19294 31950 19346
rect 32002 19294 32004 19346
rect 31948 19236 32004 19294
rect 32508 19236 32564 22652
rect 32620 22484 32676 24556
rect 32956 24052 33012 24062
rect 32956 23958 33012 23996
rect 32620 22482 33124 22484
rect 32620 22430 32622 22482
rect 32674 22430 33124 22482
rect 32620 22428 33124 22430
rect 32620 22418 32676 22428
rect 33068 22370 33124 22428
rect 33068 22318 33070 22370
rect 33122 22318 33124 22370
rect 33068 22306 33124 22318
rect 32844 22260 32900 22270
rect 32732 22258 32900 22260
rect 32732 22206 32846 22258
rect 32898 22206 32900 22258
rect 32732 22204 32900 22206
rect 32620 21812 32676 21822
rect 32732 21812 32788 22204
rect 32844 22194 32900 22204
rect 32620 21810 32788 21812
rect 32620 21758 32622 21810
rect 32674 21758 32788 21810
rect 32620 21756 32788 21758
rect 32620 21746 32676 21756
rect 33068 21700 33124 21710
rect 33068 21606 33124 21644
rect 32844 20916 32900 20926
rect 33180 20916 33236 27468
rect 33292 27076 33348 27086
rect 33404 27076 33460 27804
rect 33628 27860 33684 27870
rect 33628 27858 33908 27860
rect 33628 27806 33630 27858
rect 33682 27806 33908 27858
rect 33628 27804 33908 27806
rect 33628 27794 33684 27804
rect 33292 27074 33460 27076
rect 33292 27022 33294 27074
rect 33346 27022 33460 27074
rect 33292 27020 33460 27022
rect 33516 27748 33572 27758
rect 33292 27010 33348 27020
rect 33516 26962 33572 27692
rect 33516 26910 33518 26962
rect 33570 26910 33572 26962
rect 33516 26898 33572 26910
rect 33852 26962 33908 27804
rect 34076 27074 34132 28364
rect 34972 27860 35028 29374
rect 35644 29428 35700 29438
rect 35644 29426 35812 29428
rect 35644 29374 35646 29426
rect 35698 29374 35812 29426
rect 35644 29372 35812 29374
rect 35644 29362 35700 29372
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35756 27860 35812 29372
rect 35868 28082 35924 29708
rect 35868 28030 35870 28082
rect 35922 28030 35924 28082
rect 35868 28018 35924 28030
rect 36876 29764 36932 29774
rect 36876 28082 36932 29708
rect 36988 28644 37044 28654
rect 36988 28550 37044 28588
rect 36876 28030 36878 28082
rect 36930 28030 36932 28082
rect 36876 28018 36932 28030
rect 37324 28418 37380 31892
rect 38220 31666 38276 31892
rect 38220 31614 38222 31666
rect 38274 31614 38276 31666
rect 38220 31602 38276 31614
rect 38668 30994 38724 31006
rect 38668 30942 38670 30994
rect 38722 30942 38724 30994
rect 38108 29764 38164 29774
rect 38668 29764 38724 30942
rect 38780 30436 38836 32060
rect 38892 31108 38948 31118
rect 38892 31106 39060 31108
rect 38892 31054 38894 31106
rect 38946 31054 39060 31106
rect 38892 31052 39060 31054
rect 38892 31042 38948 31052
rect 38892 30436 38948 30446
rect 38780 30434 38948 30436
rect 38780 30382 38894 30434
rect 38946 30382 38948 30434
rect 38780 30380 38948 30382
rect 38892 30370 38948 30380
rect 38164 29708 38724 29764
rect 38108 29650 38164 29708
rect 38108 29598 38110 29650
rect 38162 29598 38164 29650
rect 38108 29586 38164 29598
rect 38892 29428 38948 29438
rect 37324 28366 37326 28418
rect 37378 28366 37380 28418
rect 36652 27860 36708 27870
rect 35756 27858 36708 27860
rect 35756 27806 36654 27858
rect 36706 27806 36708 27858
rect 35756 27804 36708 27806
rect 34972 27794 35028 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34076 27022 34078 27074
rect 34130 27022 34132 27074
rect 34076 27010 34132 27022
rect 33852 26910 33854 26962
rect 33906 26910 33908 26962
rect 33852 26898 33908 26910
rect 36540 26516 36596 27804
rect 36652 27794 36708 27804
rect 37212 27860 37268 27870
rect 37324 27860 37380 28366
rect 38556 29372 38892 29428
rect 38556 28642 38612 29372
rect 38892 29334 38948 29372
rect 39004 29316 39060 31052
rect 39116 29986 39172 29998
rect 39116 29934 39118 29986
rect 39170 29934 39172 29986
rect 39116 29652 39172 29934
rect 39564 29652 39620 29662
rect 39116 29650 39620 29652
rect 39116 29598 39118 29650
rect 39170 29598 39566 29650
rect 39618 29598 39620 29650
rect 39116 29596 39620 29598
rect 39116 29586 39172 29596
rect 39564 29586 39620 29596
rect 39676 29316 39732 32508
rect 39788 32498 39844 32508
rect 40124 32002 40180 32732
rect 40124 31950 40126 32002
rect 40178 31950 40180 32002
rect 40124 31938 40180 31950
rect 41692 32564 41748 32574
rect 41916 32564 41972 33070
rect 41692 32562 41972 32564
rect 41692 32510 41694 32562
rect 41746 32510 41972 32562
rect 41692 32508 41972 32510
rect 42252 32562 42308 33292
rect 42924 33234 42980 33292
rect 43036 33348 43092 33358
rect 43148 33348 43204 34078
rect 43484 34130 43540 34142
rect 43484 34078 43486 34130
rect 43538 34078 43540 34130
rect 43484 34020 43540 34078
rect 44156 34132 44212 34972
rect 44380 34356 44436 36428
rect 45836 36482 45892 36494
rect 45836 36430 45838 36482
rect 45890 36430 45892 36482
rect 45836 36372 45892 36430
rect 46844 36482 46900 36494
rect 46844 36430 46846 36482
rect 46898 36430 46900 36482
rect 45836 36306 45892 36316
rect 46508 36370 46564 36382
rect 46508 36318 46510 36370
rect 46562 36318 46564 36370
rect 44828 36260 44884 36270
rect 44492 36258 44884 36260
rect 44492 36206 44830 36258
rect 44882 36206 44884 36258
rect 44492 36204 44884 36206
rect 44492 35810 44548 36204
rect 44828 36194 44884 36204
rect 45164 36260 45220 36270
rect 45164 36258 45444 36260
rect 45164 36206 45166 36258
rect 45218 36206 45444 36258
rect 45164 36204 45444 36206
rect 45164 36194 45220 36204
rect 44492 35758 44494 35810
rect 44546 35758 44548 35810
rect 44492 35746 44548 35758
rect 45388 34916 45444 36204
rect 46508 35698 46564 36318
rect 46844 36372 46900 36430
rect 46844 36306 46900 36316
rect 55580 36482 55636 36494
rect 55580 36430 55582 36482
rect 55634 36430 55636 36482
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 46732 35812 46788 35822
rect 46732 35718 46788 35756
rect 55580 35812 55636 36430
rect 55580 35746 55636 35756
rect 57820 36372 57876 36382
rect 46508 35646 46510 35698
rect 46562 35646 46564 35698
rect 46508 35634 46564 35646
rect 57820 35026 57876 36316
rect 57932 35700 57988 36542
rect 57932 35634 57988 35644
rect 57820 34974 57822 35026
rect 57874 34974 57876 35026
rect 57820 34962 57876 34974
rect 45388 34850 45444 34860
rect 55580 34916 55636 34926
rect 55580 34822 55636 34860
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 44492 34356 44548 34366
rect 44380 34354 44548 34356
rect 44380 34302 44494 34354
rect 44546 34302 44548 34354
rect 44380 34300 44548 34302
rect 44492 34290 44548 34300
rect 58156 34242 58212 34254
rect 58156 34190 58158 34242
rect 58210 34190 58212 34242
rect 44156 34038 44212 34076
rect 44604 34130 44660 34142
rect 44604 34078 44606 34130
rect 44658 34078 44660 34130
rect 43484 33954 43540 33964
rect 44604 34020 44660 34078
rect 45388 34132 45444 34142
rect 44604 33954 44660 33964
rect 45276 34020 45332 34030
rect 43036 33346 43204 33348
rect 43036 33294 43038 33346
rect 43090 33294 43204 33346
rect 43036 33292 43204 33294
rect 45052 33348 45108 33358
rect 43036 33282 43092 33292
rect 45052 33254 45108 33292
rect 42924 33182 42926 33234
rect 42978 33182 42980 33234
rect 42924 33170 42980 33182
rect 42700 33124 42756 33134
rect 42252 32510 42254 32562
rect 42306 32510 42308 32562
rect 41692 30994 41748 32508
rect 42252 32498 42308 32510
rect 42364 33122 42756 33124
rect 42364 33070 42702 33122
rect 42754 33070 42756 33122
rect 42364 33068 42756 33070
rect 41692 30942 41694 30994
rect 41746 30942 41748 30994
rect 41692 30930 41748 30942
rect 41916 31108 41972 31118
rect 41916 30100 41972 31052
rect 42252 30996 42308 31006
rect 42364 30996 42420 33068
rect 42700 33058 42756 33068
rect 44828 33122 44884 33134
rect 44828 33070 44830 33122
rect 44882 33070 44884 33122
rect 44604 32676 44660 32686
rect 44828 32676 44884 33070
rect 44604 32674 44884 32676
rect 44604 32622 44606 32674
rect 44658 32622 44884 32674
rect 44604 32620 44884 32622
rect 44604 31218 44660 32620
rect 44604 31166 44606 31218
rect 44658 31166 44660 31218
rect 44604 31154 44660 31166
rect 45276 31218 45332 33964
rect 45388 32786 45444 34076
rect 58156 33684 58212 34190
rect 58156 33618 58212 33628
rect 58156 33122 58212 33134
rect 58156 33070 58158 33122
rect 58210 33070 58212 33122
rect 58156 33012 58212 33070
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 58156 32946 58212 32956
rect 50556 32890 50820 32900
rect 45388 32734 45390 32786
rect 45442 32734 45444 32786
rect 45388 32722 45444 32734
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 45276 31166 45278 31218
rect 45330 31166 45332 31218
rect 45276 31154 45332 31166
rect 57820 31108 57876 31118
rect 57820 31014 57876 31052
rect 42252 30994 42420 30996
rect 42252 30942 42254 30994
rect 42306 30942 42420 30994
rect 42252 30940 42420 30942
rect 58156 30994 58212 31006
rect 58156 30942 58158 30994
rect 58210 30942 58212 30994
rect 42252 30930 42308 30940
rect 57596 30884 57652 30894
rect 58156 30884 58212 30942
rect 57596 30882 58212 30884
rect 57596 30830 57598 30882
rect 57650 30830 58212 30882
rect 57596 30828 58212 30830
rect 57596 30818 57652 30828
rect 58156 30324 58212 30828
rect 58156 30258 58212 30268
rect 41916 30034 41972 30044
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 44492 29538 44548 29550
rect 44492 29486 44494 29538
rect 44546 29486 44548 29538
rect 41580 29428 41636 29438
rect 41580 29334 41636 29372
rect 42252 29428 42308 29438
rect 42252 29426 42644 29428
rect 42252 29374 42254 29426
rect 42306 29374 42644 29426
rect 42252 29372 42644 29374
rect 42252 29362 42308 29372
rect 39004 29314 39732 29316
rect 39004 29262 39678 29314
rect 39730 29262 39732 29314
rect 39004 29260 39732 29262
rect 38668 29204 38724 29214
rect 38668 29202 39060 29204
rect 38668 29150 38670 29202
rect 38722 29150 39060 29202
rect 38668 29148 39060 29150
rect 38668 29138 38724 29148
rect 38556 28590 38558 28642
rect 38610 28590 38612 28642
rect 37212 27858 37380 27860
rect 37212 27806 37214 27858
rect 37266 27806 37380 27858
rect 37212 27804 37380 27806
rect 37996 27860 38052 27870
rect 38556 27860 38612 28590
rect 37212 27076 37268 27804
rect 37212 27010 37268 27020
rect 37772 27300 37828 27310
rect 37772 26908 37828 27244
rect 37996 27074 38052 27804
rect 37996 27022 37998 27074
rect 38050 27022 38052 27074
rect 37996 27010 38052 27022
rect 38220 27858 38612 27860
rect 38220 27806 38558 27858
rect 38610 27806 38612 27858
rect 38220 27804 38612 27806
rect 37548 26852 37828 26908
rect 38220 26962 38276 27804
rect 38556 27794 38612 27804
rect 38220 26910 38222 26962
rect 38274 26910 38276 26962
rect 38220 26898 38276 26910
rect 36540 26514 36932 26516
rect 36540 26462 36542 26514
rect 36594 26462 36932 26514
rect 36540 26460 36932 26462
rect 36540 26450 36596 26460
rect 36204 26402 36260 26414
rect 36204 26350 36206 26402
rect 36258 26350 36260 26402
rect 34188 26068 34244 26078
rect 33852 25732 33908 25742
rect 33908 25676 34020 25732
rect 33852 25666 33908 25676
rect 33404 25506 33460 25518
rect 33404 25454 33406 25506
rect 33458 25454 33460 25506
rect 33404 24836 33460 25454
rect 33740 25506 33796 25518
rect 33740 25454 33742 25506
rect 33794 25454 33796 25506
rect 33740 25284 33796 25454
rect 33628 24836 33684 24846
rect 33404 24780 33628 24836
rect 33628 24742 33684 24780
rect 33292 24724 33348 24734
rect 33292 23828 33348 24668
rect 33404 23940 33460 23950
rect 33740 23940 33796 25228
rect 33404 23938 33796 23940
rect 33404 23886 33406 23938
rect 33458 23886 33796 23938
rect 33404 23884 33796 23886
rect 33852 24722 33908 24734
rect 33852 24670 33854 24722
rect 33906 24670 33908 24722
rect 33404 23874 33460 23884
rect 33292 23762 33348 23772
rect 33740 23044 33796 23054
rect 33628 22988 33740 23044
rect 33628 22484 33684 22988
rect 33740 22950 33796 22988
rect 33852 22708 33908 24670
rect 33964 24052 34020 25676
rect 34076 25620 34132 25630
rect 34076 25506 34132 25564
rect 34076 25454 34078 25506
rect 34130 25454 34132 25506
rect 34076 25442 34132 25454
rect 34188 24946 34244 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34636 25732 34692 25742
rect 35532 25732 35588 25742
rect 34692 25676 34804 25732
rect 34636 25666 34692 25676
rect 34188 24894 34190 24946
rect 34242 24894 34244 24946
rect 34188 24882 34244 24894
rect 34300 25282 34356 25294
rect 34300 25230 34302 25282
rect 34354 25230 34356 25282
rect 34300 24724 34356 25230
rect 34636 25282 34692 25294
rect 34636 25230 34638 25282
rect 34690 25230 34692 25282
rect 34636 25172 34692 25230
rect 34300 24658 34356 24668
rect 34412 25116 34692 25172
rect 34412 24834 34468 25116
rect 34412 24782 34414 24834
rect 34466 24782 34468 24834
rect 33964 23996 34132 24052
rect 33628 22418 33684 22428
rect 33740 22652 33908 22708
rect 33964 23828 34020 23838
rect 33404 21812 33460 21822
rect 33460 21756 33572 21812
rect 33404 21718 33460 21756
rect 33180 20860 33460 20916
rect 32844 20580 32900 20860
rect 33292 20690 33348 20702
rect 33292 20638 33294 20690
rect 33346 20638 33348 20690
rect 33292 20580 33348 20638
rect 32844 20578 33348 20580
rect 32844 20526 32846 20578
rect 32898 20526 33348 20578
rect 32844 20524 33348 20526
rect 32844 20514 32900 20524
rect 33292 20356 33348 20524
rect 33292 20290 33348 20300
rect 32732 19236 32788 19246
rect 31948 19234 32788 19236
rect 31948 19182 32734 19234
rect 32786 19182 32788 19234
rect 31948 19180 32788 19182
rect 32732 19170 32788 19180
rect 32956 19234 33012 19246
rect 32956 19182 32958 19234
rect 33010 19182 33012 19234
rect 32396 19010 32452 19022
rect 32396 18958 32398 19010
rect 32450 18958 32452 19010
rect 31948 18338 32004 18350
rect 31948 18286 31950 18338
rect 32002 18286 32004 18338
rect 31948 17780 32004 18286
rect 32172 18340 32228 18350
rect 32172 18226 32228 18284
rect 32172 18174 32174 18226
rect 32226 18174 32228 18226
rect 32172 18116 32228 18174
rect 32172 18050 32228 18060
rect 32004 17724 32116 17780
rect 31948 17714 32004 17724
rect 31948 17556 32004 17566
rect 31892 17554 32004 17556
rect 31892 17502 31950 17554
rect 32002 17502 32004 17554
rect 31892 17500 32004 17502
rect 31836 17462 31892 17500
rect 31948 17490 32004 17500
rect 32060 17220 32116 17724
rect 32060 17154 32116 17164
rect 32396 17108 32452 18958
rect 32508 18226 32564 18238
rect 32508 18174 32510 18226
rect 32562 18174 32564 18226
rect 32508 17668 32564 18174
rect 32956 17668 33012 19182
rect 33180 18676 33236 18686
rect 33180 18450 33236 18620
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 33180 18386 33236 18398
rect 33404 18450 33460 20860
rect 33516 20018 33572 21756
rect 33740 21700 33796 22652
rect 33740 21634 33796 21644
rect 33964 22370 34020 23772
rect 33964 22318 33966 22370
rect 34018 22318 34020 22370
rect 33852 21476 33908 21486
rect 33964 21476 34020 22318
rect 33852 21474 34020 21476
rect 33852 21422 33854 21474
rect 33906 21422 34020 21474
rect 33852 21420 34020 21422
rect 33852 21410 33908 21420
rect 34076 20916 34132 23996
rect 34188 23604 34244 23614
rect 34412 23604 34468 24782
rect 34524 24610 34580 24622
rect 34524 24558 34526 24610
rect 34578 24558 34580 24610
rect 34524 24500 34580 24558
rect 34636 24500 34692 24510
rect 34524 24498 34692 24500
rect 34524 24446 34638 24498
rect 34690 24446 34692 24498
rect 34524 24444 34692 24446
rect 34636 24434 34692 24444
rect 34748 23938 34804 25676
rect 35532 25618 35588 25676
rect 35532 25566 35534 25618
rect 35586 25566 35588 25618
rect 35532 25554 35588 25566
rect 35196 25506 35252 25518
rect 35196 25454 35198 25506
rect 35250 25454 35252 25506
rect 35196 24836 35252 25454
rect 35084 24724 35140 24734
rect 34972 24722 35140 24724
rect 34972 24670 35086 24722
rect 35138 24670 35140 24722
rect 34972 24668 35140 24670
rect 34860 24610 34916 24622
rect 34860 24558 34862 24610
rect 34914 24558 34916 24610
rect 34860 24500 34916 24558
rect 34860 24434 34916 24444
rect 34972 24498 35028 24668
rect 35084 24658 35140 24668
rect 35196 24500 35252 24780
rect 35644 24834 35700 24846
rect 35644 24782 35646 24834
rect 35698 24782 35700 24834
rect 35420 24724 35476 24734
rect 35420 24722 35588 24724
rect 35420 24670 35422 24722
rect 35474 24670 35588 24722
rect 35420 24668 35588 24670
rect 35420 24658 35476 24668
rect 34972 24446 34974 24498
rect 35026 24446 35028 24498
rect 34972 24434 35028 24446
rect 35084 24444 35252 24500
rect 34748 23886 34750 23938
rect 34802 23886 34804 23938
rect 34748 23828 34804 23886
rect 34748 23762 34804 23772
rect 34244 23548 34468 23604
rect 35084 23548 35140 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 24164 35588 24668
rect 35644 24612 35700 24782
rect 35644 24546 35700 24556
rect 35756 24500 35812 24510
rect 35756 24498 35924 24500
rect 35756 24446 35758 24498
rect 35810 24446 35924 24498
rect 35756 24444 35924 24446
rect 35756 24434 35812 24444
rect 35644 24164 35700 24174
rect 35532 24162 35700 24164
rect 35532 24110 35646 24162
rect 35698 24110 35700 24162
rect 35532 24108 35700 24110
rect 35644 24098 35700 24108
rect 35756 23940 35812 23950
rect 35756 23846 35812 23884
rect 35252 23828 35308 23838
rect 35308 23772 35476 23828
rect 35252 23762 35308 23772
rect 34188 23154 34244 23548
rect 34972 23492 35028 23502
rect 35084 23492 35252 23548
rect 34412 23380 34468 23390
rect 34412 23286 34468 23324
rect 34188 23102 34190 23154
rect 34242 23102 34244 23154
rect 34188 23090 34244 23102
rect 34300 23156 34356 23166
rect 34300 23062 34356 23100
rect 34524 23154 34580 23166
rect 34524 23102 34526 23154
rect 34578 23102 34580 23154
rect 34524 23044 34580 23102
rect 34748 23156 34804 23166
rect 34748 23154 34916 23156
rect 34748 23102 34750 23154
rect 34802 23102 34916 23154
rect 34748 23100 34916 23102
rect 34748 23090 34804 23100
rect 34524 22978 34580 22988
rect 34300 22258 34356 22270
rect 34300 22206 34302 22258
rect 34354 22206 34356 22258
rect 34300 21812 34356 22206
rect 34300 21746 34356 21756
rect 34524 22258 34580 22270
rect 34524 22206 34526 22258
rect 34578 22206 34580 22258
rect 34188 21586 34244 21598
rect 34188 21534 34190 21586
rect 34242 21534 34244 21586
rect 34188 21028 34244 21534
rect 34188 20962 34244 20972
rect 33852 20860 34132 20916
rect 33628 20804 33684 20814
rect 33628 20710 33684 20748
rect 33516 19966 33518 20018
rect 33570 19966 33572 20018
rect 33516 19954 33572 19966
rect 33740 20132 33796 20142
rect 33740 20018 33796 20076
rect 33740 19966 33742 20018
rect 33794 19966 33796 20018
rect 33740 19954 33796 19966
rect 33852 19236 33908 20860
rect 34076 20692 34132 20702
rect 33964 20244 34020 20254
rect 33964 19908 34020 20188
rect 34076 20130 34132 20636
rect 34300 20132 34356 20142
rect 34076 20078 34078 20130
rect 34130 20078 34132 20130
rect 34076 20066 34132 20078
rect 34188 20076 34300 20132
rect 33964 19852 34132 19908
rect 33404 18398 33406 18450
rect 33458 18398 33460 18450
rect 33180 18004 33236 18014
rect 32508 17612 33012 17668
rect 33068 17668 33124 17678
rect 32396 17042 32452 17052
rect 32508 17442 32564 17454
rect 32508 17390 32510 17442
rect 32562 17390 32564 17442
rect 31836 16770 31892 16782
rect 31836 16718 31838 16770
rect 31890 16718 31892 16770
rect 31836 16324 31892 16718
rect 31836 16258 31892 16268
rect 32060 15988 32116 15998
rect 32060 15426 32116 15932
rect 32060 15374 32062 15426
rect 32114 15374 32116 15426
rect 32060 15362 32116 15374
rect 32396 15540 32452 15550
rect 31836 15314 31892 15326
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31836 14980 31892 15262
rect 32172 15316 32228 15326
rect 32172 15202 32228 15260
rect 32172 15150 32174 15202
rect 32226 15150 32228 15202
rect 32172 15138 32228 15150
rect 31836 14914 31892 14924
rect 31724 13860 31780 14364
rect 31836 14756 31892 14766
rect 31836 13972 31892 14700
rect 31948 14644 32004 14654
rect 31948 14530 32004 14588
rect 31948 14478 31950 14530
rect 32002 14478 32004 14530
rect 31948 14466 32004 14478
rect 31836 13916 32004 13972
rect 31612 13804 31780 13860
rect 31612 12178 31668 13804
rect 31724 13636 31780 13646
rect 31724 13542 31780 13580
rect 31948 13076 32004 13916
rect 32172 13746 32228 13758
rect 32172 13694 32174 13746
rect 32226 13694 32228 13746
rect 32172 13636 32228 13694
rect 32284 13636 32340 13646
rect 32172 13580 32284 13636
rect 32284 13570 32340 13580
rect 31948 12982 32004 13020
rect 32172 12962 32228 12974
rect 32172 12910 32174 12962
rect 32226 12910 32228 12962
rect 31612 12126 31614 12178
rect 31666 12126 31668 12178
rect 31612 10948 31668 12126
rect 31724 12292 31780 12302
rect 31724 11394 31780 12236
rect 31724 11342 31726 11394
rect 31778 11342 31780 11394
rect 31724 11284 31780 11342
rect 31836 11954 31892 11966
rect 31836 11902 31838 11954
rect 31890 11902 31892 11954
rect 31836 11396 31892 11902
rect 32172 11620 32228 12910
rect 32396 12964 32452 15484
rect 32508 14532 32564 17390
rect 32620 17444 32676 17454
rect 32620 17106 32676 17388
rect 32620 17054 32622 17106
rect 32674 17054 32676 17106
rect 32620 17042 32676 17054
rect 32732 15148 32788 17612
rect 32956 17444 33012 17454
rect 32956 17350 33012 17388
rect 33068 17106 33124 17612
rect 33068 17054 33070 17106
rect 33122 17054 33124 17106
rect 33068 17042 33124 17054
rect 33180 17666 33236 17948
rect 33180 17614 33182 17666
rect 33234 17614 33236 17666
rect 33180 16996 33236 17614
rect 33180 16930 33236 16940
rect 33292 17556 33348 17566
rect 32956 16436 33012 16446
rect 32956 16210 33012 16380
rect 32956 16158 32958 16210
rect 33010 16158 33012 16210
rect 32956 16146 33012 16158
rect 33180 15316 33236 15326
rect 33180 15222 33236 15260
rect 33292 15148 33348 17500
rect 33404 17444 33460 18398
rect 33628 19234 33908 19236
rect 33628 19182 33854 19234
rect 33906 19182 33908 19234
rect 33628 19180 33908 19182
rect 33628 17668 33684 19180
rect 33852 19170 33908 19180
rect 33852 18228 33908 18238
rect 33852 18134 33908 18172
rect 33740 17780 33796 17790
rect 33740 17686 33796 17724
rect 33404 17378 33460 17388
rect 33516 17612 33684 17668
rect 33516 17220 33572 17612
rect 33628 17444 33684 17454
rect 33628 17350 33684 17388
rect 33852 17442 33908 17454
rect 33852 17390 33854 17442
rect 33906 17390 33908 17442
rect 33516 17164 33684 17220
rect 33404 17108 33460 17118
rect 33460 17052 33572 17108
rect 33404 17014 33460 17052
rect 33404 16100 33460 16110
rect 33404 16006 33460 16044
rect 33516 15148 33572 17052
rect 33628 15538 33684 17164
rect 33740 16436 33796 16446
rect 33740 16098 33796 16380
rect 33740 16046 33742 16098
rect 33794 16046 33796 16098
rect 33740 16034 33796 16046
rect 33628 15486 33630 15538
rect 33682 15486 33684 15538
rect 33628 15316 33684 15486
rect 33852 15540 33908 17390
rect 34076 16996 34132 19852
rect 34188 19012 34244 20076
rect 34300 20066 34356 20076
rect 34412 20020 34468 20030
rect 34300 19236 34356 19246
rect 34300 19142 34356 19180
rect 34412 19234 34468 19964
rect 34412 19182 34414 19234
rect 34466 19182 34468 19234
rect 34412 19170 34468 19182
rect 34188 18956 34468 19012
rect 34412 18564 34468 18956
rect 34524 18900 34580 22206
rect 34860 21812 34916 23100
rect 34972 22370 35028 23436
rect 35196 23044 35252 23492
rect 35420 23492 35476 23772
rect 35420 23378 35476 23436
rect 35420 23326 35422 23378
rect 35474 23326 35476 23378
rect 35420 23314 35476 23326
rect 35644 23714 35700 23726
rect 35644 23662 35646 23714
rect 35698 23662 35700 23714
rect 35644 23604 35700 23662
rect 35196 22978 35252 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35644 22596 35700 23548
rect 35868 23268 35924 24444
rect 36204 24164 36260 26350
rect 36876 26402 36932 26460
rect 36876 26350 36878 26402
rect 36930 26350 36932 26402
rect 36876 26338 36932 26350
rect 36988 26066 37044 26078
rect 36988 26014 36990 26066
rect 37042 26014 37044 26066
rect 36988 25284 37044 26014
rect 37324 25284 37380 25294
rect 36988 25228 37324 25284
rect 36428 24612 36484 24622
rect 36204 24098 36260 24108
rect 36316 24498 36372 24510
rect 36316 24446 36318 24498
rect 36370 24446 36372 24498
rect 36204 23940 36260 23950
rect 36316 23940 36372 24446
rect 36260 23884 36372 23940
rect 36204 23846 36260 23884
rect 35868 23202 35924 23212
rect 36204 23492 36260 23502
rect 36204 23378 36260 23436
rect 36204 23326 36206 23378
rect 36258 23326 36260 23378
rect 36204 22708 36260 23326
rect 36204 22642 36260 22652
rect 35420 22540 35700 22596
rect 34972 22318 34974 22370
rect 35026 22318 35028 22370
rect 34972 22306 35028 22318
rect 35084 22484 35140 22494
rect 34972 21812 35028 21822
rect 34860 21810 35028 21812
rect 34860 21758 34974 21810
rect 35026 21758 35028 21810
rect 34860 21756 35028 21758
rect 34972 21746 35028 21756
rect 34748 21700 34804 21710
rect 34748 21606 34804 21644
rect 34636 21586 34692 21598
rect 34636 21534 34638 21586
rect 34690 21534 34692 21586
rect 34636 20132 34692 21534
rect 35084 20916 35140 22428
rect 35308 22372 35364 22382
rect 35420 22372 35476 22540
rect 36428 22482 36484 24556
rect 36988 24610 37044 24622
rect 36988 24558 36990 24610
rect 37042 24558 37044 24610
rect 36988 24498 37044 24558
rect 36988 24446 36990 24498
rect 37042 24446 37044 24498
rect 36988 24434 37044 24446
rect 37100 24612 37156 24622
rect 36988 24164 37044 24174
rect 36764 23940 36820 23950
rect 36764 23378 36820 23884
rect 36764 23326 36766 23378
rect 36818 23326 36820 23378
rect 36764 23314 36820 23326
rect 36876 23604 36932 23614
rect 36876 23378 36932 23548
rect 36876 23326 36878 23378
rect 36930 23326 36932 23378
rect 36876 23314 36932 23326
rect 36428 22430 36430 22482
rect 36482 22430 36484 22482
rect 36428 22418 36484 22430
rect 36652 22930 36708 22942
rect 36652 22878 36654 22930
rect 36706 22878 36708 22930
rect 35308 22370 35476 22372
rect 35308 22318 35310 22370
rect 35362 22318 35476 22370
rect 35308 22316 35476 22318
rect 35308 22306 35364 22316
rect 35532 22258 35588 22270
rect 35532 22206 35534 22258
rect 35586 22206 35588 22258
rect 35420 22148 35476 22158
rect 35420 22054 35476 22092
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34636 20066 34692 20076
rect 34860 20860 35140 20916
rect 34524 18844 34692 18900
rect 34524 18676 34580 18686
rect 34524 18582 34580 18620
rect 34300 18562 34468 18564
rect 34300 18510 34414 18562
rect 34466 18510 34468 18562
rect 34300 18508 34468 18510
rect 34300 17890 34356 18508
rect 34412 18498 34468 18508
rect 34636 18116 34692 18844
rect 34860 18676 34916 20860
rect 35084 20692 35140 20702
rect 35084 20598 35140 20636
rect 35532 20468 35588 22206
rect 35980 21812 36036 21822
rect 35980 21586 36036 21756
rect 35980 21534 35982 21586
rect 36034 21534 36036 21586
rect 35980 21522 36036 21534
rect 36204 21588 36260 21598
rect 36652 21588 36708 22878
rect 36876 21700 36932 21710
rect 36876 21606 36932 21644
rect 36204 21586 36708 21588
rect 36204 21534 36206 21586
rect 36258 21534 36708 21586
rect 36204 21532 36708 21534
rect 35868 20804 35924 20814
rect 35308 20412 35588 20468
rect 35756 20748 35868 20804
rect 35196 20020 35252 20030
rect 35308 20020 35364 20412
rect 35084 20018 35364 20020
rect 35084 19966 35198 20018
rect 35250 19966 35364 20018
rect 35084 19964 35364 19966
rect 35644 20018 35700 20030
rect 35644 19966 35646 20018
rect 35698 19966 35700 20018
rect 34972 19460 35028 19470
rect 35084 19460 35140 19964
rect 35196 19954 35252 19964
rect 35420 19908 35476 19918
rect 35420 19814 35476 19852
rect 35644 19796 35700 19966
rect 35644 19730 35700 19740
rect 35756 20020 35812 20748
rect 35868 20710 35924 20748
rect 36092 20692 36148 20702
rect 36092 20598 36148 20636
rect 35868 20132 35924 20142
rect 35868 20038 35924 20076
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34972 19458 35140 19460
rect 34972 19406 34974 19458
rect 35026 19406 35140 19458
rect 34972 19404 35140 19406
rect 34972 19394 35028 19404
rect 35756 18900 35812 19964
rect 36204 20020 36260 21532
rect 36988 20916 37044 24108
rect 37100 23938 37156 24556
rect 37100 23886 37102 23938
rect 37154 23886 37156 23938
rect 37100 23604 37156 23886
rect 37100 23538 37156 23548
rect 37324 22932 37380 25228
rect 37548 23716 37604 26852
rect 38780 26740 38836 29148
rect 39004 28642 39060 29148
rect 39004 28590 39006 28642
rect 39058 28590 39060 28642
rect 39004 28578 39060 28590
rect 38892 28082 38948 28094
rect 38892 28030 38894 28082
rect 38946 28030 38948 28082
rect 38892 26962 38948 28030
rect 38892 26910 38894 26962
rect 38946 26910 38948 26962
rect 38892 26898 38948 26910
rect 39004 27858 39060 27870
rect 39004 27806 39006 27858
rect 39058 27806 39060 27858
rect 39004 26908 39060 27806
rect 39228 27860 39284 27870
rect 39228 27858 39620 27860
rect 39228 27806 39230 27858
rect 39282 27806 39620 27858
rect 39228 27804 39620 27806
rect 39228 27794 39284 27804
rect 39004 26852 39284 26908
rect 38780 26684 38948 26740
rect 37884 26572 38612 26628
rect 37884 25618 37940 26572
rect 38556 26514 38612 26572
rect 38556 26462 38558 26514
rect 38610 26462 38612 26514
rect 38556 26450 38612 26462
rect 38780 26516 38836 26526
rect 38780 26422 38836 26460
rect 37884 25566 37886 25618
rect 37938 25566 37940 25618
rect 37884 23828 37940 25566
rect 36988 20822 37044 20860
rect 37100 22876 37380 22932
rect 37436 23660 37604 23716
rect 37660 23826 37940 23828
rect 37660 23774 37886 23826
rect 37938 23774 37940 23826
rect 37660 23772 37940 23774
rect 36540 20132 36596 20142
rect 37100 20132 37156 22876
rect 37324 21588 37380 21598
rect 37212 21586 37380 21588
rect 37212 21534 37326 21586
rect 37378 21534 37380 21586
rect 37212 21532 37380 21534
rect 37212 21364 37268 21532
rect 37324 21522 37380 21532
rect 37436 21364 37492 23660
rect 37660 23266 37716 23772
rect 37884 23762 37940 23772
rect 38220 26404 38276 26414
rect 38220 26178 38276 26348
rect 38220 26126 38222 26178
rect 38274 26126 38276 26178
rect 37660 23214 37662 23266
rect 37714 23214 37716 23266
rect 37212 21298 37268 21308
rect 37324 21308 37492 21364
rect 37548 22820 37604 22830
rect 37548 21698 37604 22764
rect 37660 22036 37716 23214
rect 37772 23604 37828 23614
rect 37772 22594 37828 23548
rect 38220 23380 38276 26126
rect 38668 26178 38724 26190
rect 38668 26126 38670 26178
rect 38722 26126 38724 26178
rect 38668 26068 38724 26126
rect 38668 26002 38724 26012
rect 38780 23940 38836 23950
rect 38780 23846 38836 23884
rect 38556 23604 38612 23614
rect 38220 23324 38500 23380
rect 37996 23268 38052 23278
rect 37996 23174 38052 23212
rect 38332 23044 38388 23054
rect 38220 22930 38276 22942
rect 38220 22878 38222 22930
rect 38274 22878 38276 22930
rect 38220 22820 38276 22878
rect 38220 22754 38276 22764
rect 37772 22542 37774 22594
rect 37826 22542 37828 22594
rect 37772 22530 37828 22542
rect 38108 22484 38164 22494
rect 38108 22390 38164 22428
rect 37996 22260 38052 22270
rect 38332 22260 38388 22988
rect 37996 22258 38388 22260
rect 37996 22206 37998 22258
rect 38050 22206 38388 22258
rect 37996 22204 38388 22206
rect 37996 22194 38052 22204
rect 38444 22148 38500 23324
rect 38556 23378 38612 23548
rect 38556 23326 38558 23378
rect 38610 23326 38612 23378
rect 38556 23314 38612 23326
rect 38220 22092 38500 22148
rect 37660 21970 37716 21980
rect 38108 22036 38164 22046
rect 37548 21646 37550 21698
rect 37602 21646 37604 21698
rect 36204 19954 36260 19964
rect 36316 20018 36372 20030
rect 36316 19966 36318 20018
rect 36370 19966 36372 20018
rect 35868 19460 35924 19470
rect 35868 19346 35924 19404
rect 36316 19460 36372 19966
rect 36372 19404 36484 19460
rect 36316 19394 36372 19404
rect 35868 19294 35870 19346
rect 35922 19294 35924 19346
rect 35868 19282 35924 19294
rect 34860 18610 34916 18620
rect 35532 18844 35812 18900
rect 35196 18562 35252 18574
rect 35196 18510 35198 18562
rect 35250 18510 35252 18562
rect 34748 18452 34804 18462
rect 35084 18452 35140 18462
rect 34748 18450 35140 18452
rect 34748 18398 34750 18450
rect 34802 18398 35086 18450
rect 35138 18398 35140 18450
rect 34748 18396 35140 18398
rect 34748 18386 34804 18396
rect 35084 18386 35140 18396
rect 35196 18452 35252 18510
rect 35196 18386 35252 18396
rect 35196 18228 35252 18266
rect 35196 18162 35252 18172
rect 34636 18050 34692 18060
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17892 35588 18844
rect 35756 18676 35812 18686
rect 35756 18450 35812 18620
rect 35756 18398 35758 18450
rect 35810 18398 35812 18450
rect 35756 18386 35812 18398
rect 34300 17838 34302 17890
rect 34354 17838 34356 17890
rect 34300 17826 34356 17838
rect 35196 17836 35588 17892
rect 34524 17780 34580 17790
rect 34580 17724 34916 17780
rect 34524 17714 34580 17724
rect 34188 17554 34244 17566
rect 34188 17502 34190 17554
rect 34242 17502 34244 17554
rect 34188 17220 34244 17502
rect 34748 17556 34804 17566
rect 34748 17462 34804 17500
rect 34860 17554 34916 17724
rect 35084 17668 35140 17678
rect 35084 17574 35140 17612
rect 34860 17502 34862 17554
rect 34914 17502 34916 17554
rect 34860 17490 34916 17502
rect 34188 17154 34244 17164
rect 34300 17442 34356 17454
rect 34300 17390 34302 17442
rect 34354 17390 34356 17442
rect 34300 17108 34356 17390
rect 34300 17042 34356 17052
rect 34188 16996 34244 17006
rect 34076 16994 34244 16996
rect 34076 16942 34190 16994
rect 34242 16942 34244 16994
rect 34076 16940 34244 16942
rect 34188 16930 34244 16940
rect 34412 16996 34468 17006
rect 34412 16902 34468 16940
rect 34524 16996 34580 17006
rect 34972 16996 35028 17006
rect 34524 16994 35028 16996
rect 34524 16942 34526 16994
rect 34578 16942 34974 16994
rect 35026 16942 35028 16994
rect 34524 16940 35028 16942
rect 34524 16930 34580 16940
rect 34972 16930 35028 16940
rect 35084 16994 35140 17006
rect 35084 16942 35086 16994
rect 35138 16942 35140 16994
rect 33964 16884 34020 16894
rect 33964 16882 34132 16884
rect 33964 16830 33966 16882
rect 34018 16830 34132 16882
rect 33964 16828 34132 16830
rect 33964 16818 34020 16828
rect 34076 16436 34132 16828
rect 34412 16772 34468 16782
rect 35084 16772 35140 16942
rect 34076 16380 34356 16436
rect 34300 16210 34356 16380
rect 34300 16158 34302 16210
rect 34354 16158 34356 16210
rect 34300 16146 34356 16158
rect 33852 15484 34020 15540
rect 33740 15428 33796 15438
rect 33740 15334 33796 15372
rect 33628 15250 33684 15260
rect 33852 15314 33908 15326
rect 33852 15262 33854 15314
rect 33906 15262 33908 15314
rect 32732 15092 33124 15148
rect 33292 15092 33460 15148
rect 33516 15092 33796 15148
rect 32620 14532 32676 14542
rect 32508 14530 32676 14532
rect 32508 14478 32622 14530
rect 32674 14478 32676 14530
rect 32508 14476 32676 14478
rect 32508 13858 32564 13870
rect 32508 13806 32510 13858
rect 32562 13806 32564 13858
rect 32508 13748 32564 13806
rect 32508 13682 32564 13692
rect 32508 12964 32564 12974
rect 32396 12962 32564 12964
rect 32396 12910 32510 12962
rect 32562 12910 32564 12962
rect 32396 12908 32564 12910
rect 32172 11554 32228 11564
rect 31836 11340 32004 11396
rect 31724 11218 31780 11228
rect 31836 11172 31892 11182
rect 31836 11078 31892 11116
rect 31612 10882 31668 10892
rect 31612 10724 31668 10734
rect 31612 10630 31668 10668
rect 31500 10332 31892 10388
rect 31500 9940 31556 9950
rect 31388 9828 31444 9838
rect 31164 9826 31444 9828
rect 31164 9774 31390 9826
rect 31442 9774 31444 9826
rect 31164 9772 31444 9774
rect 31388 9762 31444 9772
rect 31500 9154 31556 9884
rect 31836 9268 31892 10332
rect 31948 9380 32004 11340
rect 32396 11394 32452 11406
rect 32396 11342 32398 11394
rect 32450 11342 32452 11394
rect 32060 11284 32116 11294
rect 32284 11284 32340 11294
rect 32060 11282 32340 11284
rect 32060 11230 32062 11282
rect 32114 11230 32286 11282
rect 32338 11230 32340 11282
rect 32060 11228 32340 11230
rect 32060 11218 32116 11228
rect 32284 11218 32340 11228
rect 32396 10834 32452 11342
rect 32396 10782 32398 10834
rect 32450 10782 32452 10834
rect 32396 10770 32452 10782
rect 32284 10610 32340 10622
rect 32284 10558 32286 10610
rect 32338 10558 32340 10610
rect 32284 10500 32340 10558
rect 32508 10500 32564 12908
rect 32284 10434 32340 10444
rect 32396 10444 32564 10500
rect 32620 10500 32676 14476
rect 32956 14420 33012 14430
rect 32732 13636 32788 13646
rect 32788 13580 32900 13636
rect 32732 13570 32788 13580
rect 31948 9324 32116 9380
rect 31500 9102 31502 9154
rect 31554 9102 31556 9154
rect 31500 9090 31556 9102
rect 31724 9212 31892 9268
rect 31052 7746 31108 7756
rect 31724 7476 31780 9212
rect 31836 9042 31892 9054
rect 31836 8990 31838 9042
rect 31890 8990 31892 9042
rect 31836 8932 31892 8990
rect 31836 8866 31892 8876
rect 30828 7474 30996 7476
rect 30828 7422 30830 7474
rect 30882 7422 30996 7474
rect 30828 7420 30996 7422
rect 31612 7474 31780 7476
rect 31612 7422 31726 7474
rect 31778 7422 31780 7474
rect 31612 7420 31780 7422
rect 30828 7410 30884 7420
rect 30716 7310 30718 7362
rect 30770 7310 30772 7362
rect 30604 7252 30660 7262
rect 30604 6578 30660 7196
rect 30604 6526 30606 6578
rect 30658 6526 30660 6578
rect 30604 6514 30660 6526
rect 30604 6020 30660 6030
rect 30604 5926 30660 5964
rect 30604 4340 30660 4350
rect 30492 4338 30660 4340
rect 30492 4286 30606 4338
rect 30658 4286 30660 4338
rect 30492 4284 30660 4286
rect 30604 4274 30660 4284
rect 29932 4228 29988 4238
rect 29708 4226 29988 4228
rect 29708 4174 29934 4226
rect 29986 4174 29988 4226
rect 29708 4172 29988 4174
rect 29932 4162 29988 4172
rect 30156 4228 30212 4238
rect 29484 3778 29652 3780
rect 29484 3726 29486 3778
rect 29538 3726 29652 3778
rect 29484 3724 29652 3726
rect 29708 3892 29764 3902
rect 29484 3714 29540 3724
rect 29036 3614 29038 3666
rect 29090 3614 29092 3666
rect 29036 3602 29092 3614
rect 28476 3490 28532 3500
rect 29708 3554 29764 3836
rect 30156 3666 30212 4172
rect 30156 3614 30158 3666
rect 30210 3614 30212 3666
rect 30156 3602 30212 3614
rect 30716 3668 30772 7310
rect 30828 6690 30884 6702
rect 30828 6638 30830 6690
rect 30882 6638 30884 6690
rect 30828 5794 30884 6638
rect 31500 6468 31556 6478
rect 31164 5908 31220 5918
rect 31500 5908 31556 6412
rect 31164 5814 31220 5852
rect 31276 5906 31556 5908
rect 31276 5854 31502 5906
rect 31554 5854 31556 5906
rect 31276 5852 31556 5854
rect 30828 5742 30830 5794
rect 30882 5742 30884 5794
rect 30828 5730 30884 5742
rect 31276 5460 31332 5852
rect 31500 5842 31556 5852
rect 30828 5122 30884 5134
rect 30828 5070 30830 5122
rect 30882 5070 30884 5122
rect 30828 3892 30884 5070
rect 30940 4788 30996 4798
rect 30940 4450 30996 4732
rect 30940 4398 30942 4450
rect 30994 4398 30996 4450
rect 30940 4386 30996 4398
rect 30828 3826 30884 3836
rect 30828 3668 30884 3678
rect 30716 3666 30884 3668
rect 30716 3614 30830 3666
rect 30882 3614 30884 3666
rect 30716 3612 30884 3614
rect 30828 3602 30884 3612
rect 31276 3666 31332 5404
rect 31500 5348 31556 5358
rect 31500 4338 31556 5292
rect 31612 5346 31668 7420
rect 31724 7410 31780 7420
rect 31836 8484 31892 8494
rect 31612 5294 31614 5346
rect 31666 5294 31668 5346
rect 31612 5236 31668 5294
rect 31612 5170 31668 5180
rect 31724 5796 31780 5806
rect 31612 4564 31668 4574
rect 31724 4564 31780 5740
rect 31836 5684 31892 8428
rect 31948 8146 32004 8158
rect 31948 8094 31950 8146
rect 32002 8094 32004 8146
rect 31948 7250 32004 8094
rect 31948 7198 31950 7250
rect 32002 7198 32004 7250
rect 31948 7186 32004 7198
rect 32060 6580 32116 9324
rect 32396 9156 32452 10444
rect 32620 10434 32676 10444
rect 32732 12740 32788 12750
rect 32508 10276 32564 10286
rect 32508 9826 32564 10220
rect 32508 9774 32510 9826
rect 32562 9774 32564 9826
rect 32508 9762 32564 9774
rect 32396 9090 32452 9100
rect 32396 8260 32452 8270
rect 32396 8258 32564 8260
rect 32396 8206 32398 8258
rect 32450 8206 32564 8258
rect 32396 8204 32564 8206
rect 32396 8194 32452 8204
rect 32508 8036 32564 8204
rect 32284 7476 32340 7486
rect 32284 7474 32452 7476
rect 32284 7422 32286 7474
rect 32338 7422 32452 7474
rect 32284 7420 32452 7422
rect 32284 7410 32340 7420
rect 32284 6692 32340 6702
rect 32284 6598 32340 6636
rect 32172 6580 32228 6590
rect 32060 6524 32172 6580
rect 32172 6514 32228 6524
rect 32172 6020 32228 6030
rect 31948 5908 32004 5918
rect 31948 5814 32004 5852
rect 32172 5684 32228 5964
rect 31836 5618 31892 5628
rect 31948 5628 32228 5684
rect 32284 5908 32340 5918
rect 32396 5908 32452 7420
rect 32284 5906 32452 5908
rect 32284 5854 32286 5906
rect 32338 5854 32452 5906
rect 32284 5852 32452 5854
rect 31612 4562 31780 4564
rect 31612 4510 31614 4562
rect 31666 4510 31780 4562
rect 31612 4508 31780 4510
rect 31612 4498 31668 4508
rect 31500 4286 31502 4338
rect 31554 4286 31556 4338
rect 31500 4274 31556 4286
rect 31948 4228 32004 5628
rect 32060 5348 32116 5358
rect 32060 5234 32116 5292
rect 32060 5182 32062 5234
rect 32114 5182 32116 5234
rect 32060 5170 32116 5182
rect 32172 5122 32228 5134
rect 32172 5070 32174 5122
rect 32226 5070 32228 5122
rect 32172 5012 32228 5070
rect 32284 5124 32340 5852
rect 32396 5124 32452 5134
rect 32284 5068 32396 5124
rect 32172 4946 32228 4956
rect 32172 4228 32228 4238
rect 31948 4172 32172 4228
rect 32172 4134 32228 4172
rect 31276 3614 31278 3666
rect 31330 3614 31332 3666
rect 31276 3602 31332 3614
rect 29708 3502 29710 3554
rect 29762 3502 29764 3554
rect 29708 3490 29764 3502
rect 31612 3556 31668 3566
rect 29484 3444 29540 3482
rect 31612 3462 31668 3500
rect 29484 2884 29540 3388
rect 32396 3444 32452 5068
rect 32396 3378 32452 3388
rect 29484 2818 29540 2828
rect 32508 2436 32564 7980
rect 32620 6020 32676 6030
rect 32732 6020 32788 12684
rect 32844 7476 32900 13580
rect 32956 13186 33012 14364
rect 32956 13134 32958 13186
rect 33010 13134 33012 13186
rect 32956 13122 33012 13134
rect 33068 12290 33124 15092
rect 33292 14754 33348 14766
rect 33292 14702 33294 14754
rect 33346 14702 33348 14754
rect 33180 13636 33236 13646
rect 33180 13542 33236 13580
rect 33292 12404 33348 14702
rect 33404 13412 33460 15092
rect 33404 13346 33460 13356
rect 33516 14980 33572 14990
rect 33516 12850 33572 14924
rect 33628 14530 33684 14542
rect 33628 14478 33630 14530
rect 33682 14478 33684 14530
rect 33628 13300 33684 14478
rect 33740 14420 33796 15092
rect 33852 14642 33908 15262
rect 33964 15204 34020 15484
rect 34076 15428 34132 15438
rect 34300 15428 34356 15438
rect 34132 15426 34356 15428
rect 34132 15374 34302 15426
rect 34354 15374 34356 15426
rect 34132 15372 34356 15374
rect 34076 15362 34132 15372
rect 34300 15362 34356 15372
rect 34412 15426 34468 16716
rect 34636 16716 35140 16772
rect 34636 15538 34692 16716
rect 35196 16660 35252 17836
rect 36428 17780 36484 19404
rect 36540 19012 36596 20076
rect 36764 20076 37156 20132
rect 37212 20802 37268 20814
rect 37212 20750 37214 20802
rect 37266 20750 37268 20802
rect 36764 19684 36820 20076
rect 36876 19908 36932 19918
rect 36876 19796 36932 19852
rect 37100 19796 37156 19806
rect 36876 19794 37156 19796
rect 36876 19742 37102 19794
rect 37154 19742 37156 19794
rect 36876 19740 37156 19742
rect 37100 19730 37156 19740
rect 37212 19796 37268 20750
rect 36764 19628 37044 19684
rect 36540 18946 36596 18956
rect 36652 17892 36708 17902
rect 36540 17780 36596 17790
rect 36428 17724 36540 17780
rect 36540 17686 36596 17724
rect 35980 17442 36036 17454
rect 35980 17390 35982 17442
rect 36034 17390 36036 17442
rect 35980 17332 36036 17390
rect 35980 17266 36036 17276
rect 35308 16882 35364 16894
rect 35308 16830 35310 16882
rect 35362 16830 35364 16882
rect 35308 16772 35364 16830
rect 35308 16706 35364 16716
rect 35196 16594 35252 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 36540 15874 36596 15886
rect 36540 15822 36542 15874
rect 36594 15822 36596 15874
rect 34636 15486 34638 15538
rect 34690 15486 34692 15538
rect 34636 15474 34692 15486
rect 35868 15652 35924 15662
rect 35868 15538 35924 15596
rect 35868 15486 35870 15538
rect 35922 15486 35924 15538
rect 35868 15474 35924 15486
rect 34412 15374 34414 15426
rect 34466 15374 34468 15426
rect 33964 15148 34132 15204
rect 33852 14590 33854 14642
rect 33906 14590 33908 14642
rect 33852 14578 33908 14590
rect 33964 14530 34020 14542
rect 33964 14478 33966 14530
rect 34018 14478 34020 14530
rect 33964 14420 34020 14478
rect 34076 14532 34132 15148
rect 34412 15092 34468 15374
rect 36428 15426 36484 15438
rect 36428 15374 36430 15426
rect 36482 15374 36484 15426
rect 34412 15026 34468 15036
rect 34636 15316 34692 15326
rect 34188 14532 34244 14542
rect 34076 14530 34244 14532
rect 34076 14478 34190 14530
rect 34242 14478 34244 14530
rect 34076 14476 34244 14478
rect 33740 14364 34020 14420
rect 34188 14420 34244 14476
rect 33628 13234 33684 13244
rect 33740 13746 33796 13758
rect 33740 13694 33742 13746
rect 33794 13694 33796 13746
rect 33740 13074 33796 13694
rect 33852 13524 33908 14364
rect 34188 14354 34244 14364
rect 34636 14418 34692 15260
rect 34972 15314 35028 15326
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34972 15148 35028 15262
rect 36092 15314 36148 15326
rect 36092 15262 36094 15314
rect 36146 15262 36148 15314
rect 34972 15092 35140 15148
rect 34972 15026 35028 15036
rect 34636 14366 34638 14418
rect 34690 14366 34692 14418
rect 34636 14354 34692 14366
rect 34748 14308 34804 14318
rect 33852 13458 33908 13468
rect 34076 13860 34132 13870
rect 33740 13022 33742 13074
rect 33794 13022 33796 13074
rect 33740 13010 33796 13022
rect 33516 12798 33518 12850
rect 33570 12798 33572 12850
rect 33516 12740 33572 12798
rect 33516 12674 33572 12684
rect 33964 12962 34020 12974
rect 33964 12910 33966 12962
rect 34018 12910 34020 12962
rect 33964 12740 34020 12910
rect 33964 12674 34020 12684
rect 33292 12348 33572 12404
rect 33068 12238 33070 12290
rect 33122 12238 33124 12290
rect 33068 12226 33124 12238
rect 33292 12178 33348 12190
rect 33292 12126 33294 12178
rect 33346 12126 33348 12178
rect 33292 10724 33348 12126
rect 33292 10658 33348 10668
rect 33404 11954 33460 11966
rect 33404 11902 33406 11954
rect 33458 11902 33460 11954
rect 33404 10610 33460 11902
rect 33404 10558 33406 10610
rect 33458 10558 33460 10610
rect 33404 10546 33460 10558
rect 33404 10052 33460 10062
rect 33404 9958 33460 9996
rect 32956 9938 33012 9950
rect 32956 9886 32958 9938
rect 33010 9886 33012 9938
rect 32956 9604 33012 9886
rect 32956 8820 33012 9548
rect 33404 9716 33460 9726
rect 33180 9156 33236 9166
rect 33180 9062 33236 9100
rect 33068 9044 33124 9054
rect 33068 8950 33124 8988
rect 32956 8754 33012 8764
rect 33404 8034 33460 9660
rect 33516 8260 33572 12348
rect 34076 12290 34132 13804
rect 34748 13748 34804 14252
rect 34972 14306 35028 14318
rect 34972 14254 34974 14306
rect 35026 14254 35028 14306
rect 34972 14196 35028 14254
rect 34972 14130 35028 14140
rect 34636 13746 34804 13748
rect 34636 13694 34750 13746
rect 34802 13694 34804 13746
rect 34636 13692 34804 13694
rect 34300 13188 34356 13198
rect 34300 12962 34356 13132
rect 34300 12910 34302 12962
rect 34354 12910 34356 12962
rect 34300 12898 34356 12910
rect 34636 12404 34692 13692
rect 34748 13682 34804 13692
rect 35084 13636 35140 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 36092 14418 36148 15262
rect 36428 14756 36484 15374
rect 36092 14366 36094 14418
rect 36146 14366 36148 14418
rect 35420 14308 35476 14318
rect 35420 14214 35476 14252
rect 35532 13748 35588 13758
rect 36092 13748 36148 14366
rect 36204 14700 36428 14756
rect 36204 14418 36260 14700
rect 36428 14690 36484 14700
rect 36428 14532 36484 14542
rect 36428 14438 36484 14476
rect 36204 14366 36206 14418
rect 36258 14366 36260 14418
rect 36204 14354 36260 14366
rect 36540 14308 36596 15822
rect 36652 15148 36708 17836
rect 36876 17108 36932 17118
rect 36876 16884 36932 17052
rect 36988 16996 37044 19628
rect 37100 18900 37156 18910
rect 37212 18900 37268 19740
rect 37156 18844 37268 18900
rect 37100 17108 37156 18844
rect 37212 17666 37268 17678
rect 37212 17614 37214 17666
rect 37266 17614 37268 17666
rect 37212 17332 37268 17614
rect 37212 17266 37268 17276
rect 37100 17052 37268 17108
rect 36988 16940 37156 16996
rect 36876 16828 37044 16884
rect 36988 16770 37044 16828
rect 36988 16718 36990 16770
rect 37042 16718 37044 16770
rect 36988 16706 37044 16718
rect 37100 16548 37156 16940
rect 36988 16492 37156 16548
rect 36988 15876 37044 16492
rect 36876 15820 37044 15876
rect 37100 15876 37156 15886
rect 36876 15428 36932 15820
rect 37100 15782 37156 15820
rect 36876 15362 36932 15372
rect 36988 15652 37044 15662
rect 36988 15314 37044 15596
rect 37100 15540 37156 15550
rect 37100 15446 37156 15484
rect 36988 15262 36990 15314
rect 37042 15262 37044 15314
rect 36988 15204 37044 15262
rect 36652 15092 36820 15148
rect 36988 15138 37044 15148
rect 36652 14308 36708 14318
rect 36540 14252 36652 14308
rect 36652 14242 36708 14252
rect 36428 14196 36484 14206
rect 36484 14140 36596 14196
rect 36428 14130 36484 14140
rect 36092 13692 36260 13748
rect 35532 13654 35588 13692
rect 35084 13074 35140 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13022 35086 13074
rect 35138 13022 35140 13074
rect 35084 13010 35140 13022
rect 35868 13074 35924 13086
rect 35868 13022 35870 13074
rect 35922 13022 35924 13074
rect 35644 12964 35700 12974
rect 34076 12238 34078 12290
rect 34130 12238 34132 12290
rect 34076 12226 34132 12238
rect 34188 12348 34692 12404
rect 35532 12850 35588 12862
rect 35532 12798 35534 12850
rect 35586 12798 35588 12850
rect 34188 10724 34244 12348
rect 34524 12178 34580 12190
rect 34524 12126 34526 12178
rect 34578 12126 34580 12178
rect 34524 11620 34580 12126
rect 34524 11554 34580 11564
rect 34636 12180 34692 12190
rect 34636 11396 34692 12124
rect 35084 12180 35140 12190
rect 35084 12086 35140 12124
rect 33964 10668 34244 10724
rect 34300 11394 34692 11396
rect 34300 11342 34638 11394
rect 34690 11342 34692 11394
rect 34300 11340 34692 11342
rect 33852 10498 33908 10510
rect 33852 10446 33854 10498
rect 33906 10446 33908 10498
rect 33740 8596 33796 8606
rect 33628 8260 33684 8270
rect 33516 8258 33684 8260
rect 33516 8206 33630 8258
rect 33682 8206 33684 8258
rect 33516 8204 33684 8206
rect 33628 8194 33684 8204
rect 33404 7982 33406 8034
rect 33458 7982 33460 8034
rect 33404 7970 33460 7982
rect 33740 7812 33796 8540
rect 33852 8484 33908 10446
rect 33852 8418 33908 8428
rect 33964 7812 34020 10668
rect 34300 10612 34356 11340
rect 34524 10724 34580 10734
rect 34524 10630 34580 10668
rect 34188 10610 34356 10612
rect 34188 10558 34302 10610
rect 34354 10558 34356 10610
rect 34188 10556 34356 10558
rect 34076 9266 34132 9278
rect 34076 9214 34078 9266
rect 34130 9214 34132 9266
rect 34076 8146 34132 9214
rect 34188 9042 34244 10556
rect 34300 10546 34356 10556
rect 34636 9940 34692 11340
rect 34860 11844 34916 11854
rect 34748 9940 34804 9950
rect 34636 9938 34804 9940
rect 34636 9886 34750 9938
rect 34802 9886 34804 9938
rect 34636 9884 34804 9886
rect 34748 9874 34804 9884
rect 34300 9828 34356 9838
rect 34300 9734 34356 9772
rect 34188 8990 34190 9042
rect 34242 8990 34244 9042
rect 34188 8978 34244 8990
rect 34636 8932 34692 8942
rect 34636 8596 34692 8876
rect 34636 8530 34692 8540
rect 34076 8094 34078 8146
rect 34130 8094 34132 8146
rect 34076 8082 34132 8094
rect 33628 7756 33796 7812
rect 33852 7756 34020 7812
rect 32844 7410 32900 7420
rect 33180 7474 33236 7486
rect 33180 7422 33182 7474
rect 33234 7422 33236 7474
rect 32676 5964 32788 6020
rect 33180 6916 33236 7422
rect 32620 5954 32676 5964
rect 33180 5012 33236 6860
rect 33516 6804 33572 6814
rect 33516 5572 33572 6748
rect 33628 6244 33684 7756
rect 33740 7476 33796 7486
rect 33740 7382 33796 7420
rect 33852 6468 33908 7756
rect 34076 7476 34132 7486
rect 33852 6402 33908 6412
rect 33964 7474 34132 7476
rect 33964 7422 34078 7474
rect 34130 7422 34132 7474
rect 33964 7420 34132 7422
rect 33628 6188 33908 6244
rect 33628 6018 33684 6030
rect 33628 5966 33630 6018
rect 33682 5966 33684 6018
rect 33628 5796 33684 5966
rect 33628 5730 33684 5740
rect 33852 5684 33908 6188
rect 33964 5908 34020 7420
rect 34076 7410 34132 7420
rect 34300 7474 34356 7486
rect 34300 7422 34302 7474
rect 34354 7422 34356 7474
rect 34188 7364 34244 7374
rect 34188 7270 34244 7308
rect 34076 6690 34132 6702
rect 34076 6638 34078 6690
rect 34130 6638 34132 6690
rect 34076 6580 34132 6638
rect 34076 6514 34132 6524
rect 33964 5842 34020 5852
rect 34076 6132 34132 6142
rect 34300 6132 34356 7422
rect 34748 7476 34804 7486
rect 34860 7476 34916 11788
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34972 11620 35028 11630
rect 34972 10052 35028 11564
rect 35084 11284 35140 11294
rect 35084 10834 35140 11228
rect 35532 11172 35588 12798
rect 35644 12290 35700 12908
rect 35644 12238 35646 12290
rect 35698 12238 35700 12290
rect 35644 12226 35700 12238
rect 35756 12738 35812 12750
rect 35756 12686 35758 12738
rect 35810 12686 35812 12738
rect 35756 11620 35812 12686
rect 35868 12180 35924 13022
rect 35868 12114 35924 12124
rect 35532 11106 35588 11116
rect 35644 11564 35812 11620
rect 35868 11956 35924 11966
rect 35084 10782 35086 10834
rect 35138 10782 35140 10834
rect 35084 10770 35140 10782
rect 35644 10836 35700 11564
rect 35644 10610 35700 10780
rect 35644 10558 35646 10610
rect 35698 10558 35700 10610
rect 35644 10546 35700 10558
rect 35756 10612 35812 10622
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34972 9996 35364 10052
rect 35084 9828 35140 9838
rect 34972 8036 35028 8046
rect 34972 7942 35028 7980
rect 35084 7698 35140 9772
rect 35308 9602 35364 9996
rect 35756 9938 35812 10556
rect 35756 9886 35758 9938
rect 35810 9886 35812 9938
rect 35756 9874 35812 9886
rect 35868 9940 35924 11900
rect 36092 11508 36148 11518
rect 36204 11508 36260 13692
rect 36148 11452 36260 11508
rect 36316 12740 36372 12750
rect 36092 11442 36148 11452
rect 36316 11394 36372 12684
rect 36428 12180 36484 12190
rect 36428 12086 36484 12124
rect 36316 11342 36318 11394
rect 36370 11342 36372 11394
rect 36204 11172 36260 11182
rect 36204 10722 36260 11116
rect 36204 10670 36206 10722
rect 36258 10670 36260 10722
rect 36204 10658 36260 10670
rect 35308 9550 35310 9602
rect 35362 9550 35364 9602
rect 35308 8820 35364 9550
rect 35868 9154 35924 9884
rect 36204 9604 36260 9614
rect 36204 9510 36260 9548
rect 36316 9380 36372 11342
rect 36428 11284 36484 11294
rect 36540 11284 36596 14140
rect 36428 11282 36596 11284
rect 36428 11230 36430 11282
rect 36482 11230 36596 11282
rect 36428 11228 36596 11230
rect 36428 11218 36484 11228
rect 36764 10388 36820 15092
rect 37100 15092 37156 15102
rect 37100 14644 37156 15036
rect 36988 14588 37156 14644
rect 36988 13746 37044 14588
rect 37100 14420 37156 14430
rect 37100 14326 37156 14364
rect 36988 13694 36990 13746
rect 37042 13694 37044 13746
rect 36988 13682 37044 13694
rect 37100 13636 37156 13646
rect 37100 13542 37156 13580
rect 37100 12852 37156 12862
rect 37100 12758 37156 12796
rect 36876 12066 36932 12078
rect 36876 12014 36878 12066
rect 36930 12014 36932 12066
rect 36876 11508 36932 12014
rect 36876 11442 36932 11452
rect 37100 11394 37156 11406
rect 37100 11342 37102 11394
rect 37154 11342 37156 11394
rect 37100 10724 37156 11342
rect 37212 10834 37268 17052
rect 37324 15652 37380 21308
rect 37548 21026 37604 21646
rect 38108 21586 38164 21980
rect 38108 21534 38110 21586
rect 38162 21534 38164 21586
rect 38108 21522 38164 21534
rect 38220 21364 38276 22092
rect 37548 20974 37550 21026
rect 37602 20974 37604 21026
rect 37548 20962 37604 20974
rect 38108 21308 38276 21364
rect 38444 21364 38500 21374
rect 37996 20804 38052 20814
rect 37996 20710 38052 20748
rect 37436 20132 37492 20142
rect 37436 20038 37492 20076
rect 37996 20020 38052 20030
rect 37996 19926 38052 19964
rect 37884 19794 37940 19806
rect 37884 19742 37886 19794
rect 37938 19742 37940 19794
rect 37436 19012 37492 19022
rect 37436 16660 37492 18956
rect 37884 18900 37940 19742
rect 37884 18834 37940 18844
rect 37996 18452 38052 18462
rect 37996 18358 38052 18396
rect 37772 18116 37828 18126
rect 37660 18060 37772 18116
rect 37548 17780 37604 17790
rect 37548 17686 37604 17724
rect 37548 16884 37604 16894
rect 37548 16790 37604 16828
rect 37436 16604 37604 16660
rect 37436 15986 37492 15998
rect 37436 15934 37438 15986
rect 37490 15934 37492 15986
rect 37436 15876 37492 15934
rect 37436 15810 37492 15820
rect 37436 15652 37492 15662
rect 37324 15596 37436 15652
rect 37436 15586 37492 15596
rect 37324 15428 37380 15438
rect 37324 14756 37380 15372
rect 37548 14980 37604 16604
rect 37660 15092 37716 18060
rect 37772 18050 37828 18060
rect 37772 17554 37828 17566
rect 37772 17502 37774 17554
rect 37826 17502 37828 17554
rect 37772 16884 37828 17502
rect 37772 16818 37828 16828
rect 37884 17554 37940 17566
rect 37884 17502 37886 17554
rect 37938 17502 37940 17554
rect 37772 16324 37828 16334
rect 37884 16324 37940 17502
rect 38108 17108 38164 21308
rect 38444 21270 38500 21308
rect 38220 20916 38276 20926
rect 38444 20916 38500 20926
rect 38276 20914 38500 20916
rect 38276 20862 38446 20914
rect 38498 20862 38500 20914
rect 38276 20860 38500 20862
rect 38220 20850 38276 20860
rect 38220 20018 38276 20030
rect 38220 19966 38222 20018
rect 38274 19966 38276 20018
rect 38220 19012 38276 19966
rect 38444 19684 38500 20860
rect 38444 19618 38500 19628
rect 38220 18946 38276 18956
rect 38332 18452 38388 18462
rect 38668 18452 38724 18462
rect 38892 18452 38948 26684
rect 39228 26516 39284 26852
rect 39116 26460 39284 26516
rect 39564 26514 39620 27804
rect 39676 26628 39732 29260
rect 42588 28642 42644 29372
rect 42588 28590 42590 28642
rect 42642 28590 42644 28642
rect 42588 28578 42644 28590
rect 43372 29204 43428 29214
rect 41020 28532 41076 28542
rect 39676 26562 39732 26572
rect 40236 27188 40292 27198
rect 39564 26462 39566 26514
rect 39618 26462 39620 26514
rect 39004 25508 39060 25518
rect 39004 25414 39060 25452
rect 39116 23156 39172 26460
rect 39564 26450 39620 26462
rect 40236 26514 40292 27132
rect 41020 27188 41076 28476
rect 41580 28532 41636 28542
rect 41580 28418 41636 28476
rect 42924 28532 42980 28542
rect 43148 28532 43204 28542
rect 42924 28530 43204 28532
rect 42924 28478 42926 28530
rect 42978 28478 43150 28530
rect 43202 28478 43204 28530
rect 42924 28476 43204 28478
rect 42924 28466 42980 28476
rect 43148 28466 43204 28476
rect 43372 28530 43428 29148
rect 43932 28644 43988 28654
rect 43596 28642 43988 28644
rect 43596 28590 43934 28642
rect 43986 28590 43988 28642
rect 43596 28588 43988 28590
rect 43372 28478 43374 28530
rect 43426 28478 43428 28530
rect 41580 28366 41582 28418
rect 41634 28366 41636 28418
rect 41580 28354 41636 28366
rect 42028 28420 42084 28430
rect 41356 27860 41412 27870
rect 41356 27766 41412 27804
rect 42028 27858 42084 28364
rect 42140 28420 42196 28430
rect 42812 28420 42868 28430
rect 42140 28418 42420 28420
rect 42140 28366 42142 28418
rect 42194 28366 42420 28418
rect 42140 28364 42420 28366
rect 42140 28354 42196 28364
rect 42028 27806 42030 27858
rect 42082 27806 42084 27858
rect 42028 27794 42084 27806
rect 42252 27636 42308 27646
rect 41020 27094 41076 27132
rect 42140 27580 42252 27636
rect 41468 27076 41524 27086
rect 41468 26982 41524 27020
rect 40684 26852 40740 26862
rect 40236 26462 40238 26514
rect 40290 26462 40292 26514
rect 40236 26450 40292 26462
rect 40348 26850 40740 26852
rect 40348 26798 40686 26850
rect 40738 26798 40740 26850
rect 40348 26796 40740 26798
rect 39676 26404 39732 26414
rect 39676 26310 39732 26348
rect 40348 26402 40404 26796
rect 40684 26786 40740 26796
rect 42140 26516 42196 27580
rect 42252 27570 42308 27580
rect 40348 26350 40350 26402
rect 40402 26350 40404 26402
rect 40348 26338 40404 26350
rect 41916 26514 42196 26516
rect 41916 26462 42142 26514
rect 42194 26462 42196 26514
rect 41916 26460 42196 26462
rect 39228 26292 39284 26302
rect 39228 26290 39620 26292
rect 39228 26238 39230 26290
rect 39282 26238 39620 26290
rect 39228 26236 39620 26238
rect 39228 26226 39284 26236
rect 39564 26180 39620 26236
rect 40012 26290 40068 26302
rect 40012 26238 40014 26290
rect 40066 26238 40068 26290
rect 40012 26180 40068 26238
rect 39564 26124 40068 26180
rect 39228 26068 39284 26078
rect 39452 26068 39508 26078
rect 39284 26066 39508 26068
rect 39284 26014 39454 26066
rect 39506 26014 39508 26066
rect 39284 26012 39508 26014
rect 39228 26002 39284 26012
rect 39452 26002 39508 26012
rect 39564 25506 39620 26124
rect 39564 25454 39566 25506
rect 39618 25454 39620 25506
rect 39564 25442 39620 25454
rect 40236 25394 40292 25406
rect 40236 25342 40238 25394
rect 40290 25342 40292 25394
rect 40236 23604 40292 25342
rect 41244 25284 41300 25294
rect 40796 23938 40852 23950
rect 40796 23886 40798 23938
rect 40850 23886 40852 23938
rect 40348 23828 40404 23838
rect 40348 23734 40404 23772
rect 40236 23548 40404 23604
rect 40012 23268 40068 23278
rect 39116 23100 39620 23156
rect 39004 23044 39060 23054
rect 39004 22950 39060 22988
rect 39116 22932 39172 22942
rect 39004 22708 39060 22718
rect 39004 22482 39060 22652
rect 39116 22596 39172 22876
rect 39228 22930 39284 22942
rect 39228 22878 39230 22930
rect 39282 22878 39284 22930
rect 39228 22820 39284 22878
rect 39228 22754 39284 22764
rect 39452 22930 39508 22942
rect 39452 22878 39454 22930
rect 39506 22878 39508 22930
rect 39228 22596 39284 22606
rect 39116 22594 39284 22596
rect 39116 22542 39230 22594
rect 39282 22542 39284 22594
rect 39116 22540 39284 22542
rect 39228 22530 39284 22540
rect 39004 22430 39006 22482
rect 39058 22430 39060 22482
rect 39004 22418 39060 22430
rect 39452 22370 39508 22878
rect 39452 22318 39454 22370
rect 39506 22318 39508 22370
rect 39452 21924 39508 22318
rect 39452 21858 39508 21868
rect 38332 18450 38948 18452
rect 38332 18398 38334 18450
rect 38386 18398 38670 18450
rect 38722 18398 38948 18450
rect 38332 18396 38948 18398
rect 39564 18674 39620 23100
rect 39676 22932 39732 22942
rect 39676 22838 39732 22876
rect 39788 22708 39844 22718
rect 39788 22370 39844 22652
rect 40012 22482 40068 23212
rect 40124 23156 40180 23166
rect 40124 23062 40180 23100
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 40012 22418 40068 22430
rect 40124 22820 40180 22830
rect 39788 22318 39790 22370
rect 39842 22318 39844 22370
rect 39788 22306 39844 22318
rect 40124 22370 40180 22764
rect 40124 22318 40126 22370
rect 40178 22318 40180 22370
rect 40124 22306 40180 22318
rect 39900 22146 39956 22158
rect 39900 22094 39902 22146
rect 39954 22094 39956 22146
rect 39900 20914 39956 22094
rect 39900 20862 39902 20914
rect 39954 20862 39956 20914
rect 39900 20850 39956 20862
rect 40012 20692 40068 20702
rect 40236 20692 40292 20702
rect 40012 20690 40292 20692
rect 40012 20638 40014 20690
rect 40066 20638 40238 20690
rect 40290 20638 40292 20690
rect 40012 20636 40292 20638
rect 40012 20626 40068 20636
rect 40236 20626 40292 20636
rect 39788 20580 39844 20590
rect 39564 18622 39566 18674
rect 39618 18622 39620 18674
rect 38332 18386 38388 18396
rect 38668 18358 38724 18396
rect 39228 18340 39284 18350
rect 39564 18340 39620 18622
rect 39228 18338 39396 18340
rect 39228 18286 39230 18338
rect 39282 18286 39396 18338
rect 39228 18284 39396 18286
rect 39228 18274 39284 18284
rect 38444 18228 38500 18238
rect 38500 18172 38612 18228
rect 38444 18162 38500 18172
rect 38220 17556 38276 17566
rect 38444 17556 38500 17566
rect 38220 17554 38500 17556
rect 38220 17502 38222 17554
rect 38274 17502 38446 17554
rect 38498 17502 38500 17554
rect 38220 17500 38500 17502
rect 38220 17490 38276 17500
rect 38444 17490 38500 17500
rect 38108 17042 38164 17052
rect 37772 16322 37940 16324
rect 37772 16270 37774 16322
rect 37826 16270 37940 16322
rect 37772 16268 37940 16270
rect 37996 16996 38052 17006
rect 37772 16258 37828 16268
rect 37996 16212 38052 16940
rect 37884 16156 38052 16212
rect 38220 16994 38276 17006
rect 38220 16942 38222 16994
rect 38274 16942 38276 16994
rect 37772 16100 37828 16110
rect 37884 16100 37940 16156
rect 38220 16100 38276 16942
rect 37772 16098 37940 16100
rect 37772 16046 37774 16098
rect 37826 16046 37940 16098
rect 37772 16044 37940 16046
rect 37996 16044 38276 16100
rect 38332 16882 38388 16894
rect 38332 16830 38334 16882
rect 38386 16830 38388 16882
rect 37772 16034 37828 16044
rect 37884 15876 37940 15886
rect 37884 15538 37940 15820
rect 37884 15486 37886 15538
rect 37938 15486 37940 15538
rect 37884 15474 37940 15486
rect 37660 15026 37716 15036
rect 37548 14914 37604 14924
rect 37324 14700 37940 14756
rect 37884 14532 37940 14700
rect 37996 14754 38052 16044
rect 38220 15876 38276 15886
rect 38108 15652 38164 15662
rect 38108 15148 38164 15596
rect 38220 15314 38276 15820
rect 38332 15540 38388 16830
rect 38556 15988 38612 18172
rect 38780 17668 38836 17678
rect 39340 17668 39396 18284
rect 38780 17574 38836 17612
rect 39228 17666 39396 17668
rect 39228 17614 39342 17666
rect 39394 17614 39396 17666
rect 39228 17612 39396 17614
rect 39004 17554 39060 17566
rect 39004 17502 39006 17554
rect 39058 17502 39060 17554
rect 38892 17442 38948 17454
rect 38892 17390 38894 17442
rect 38946 17390 38948 17442
rect 38892 17332 38948 17390
rect 38892 17266 38948 17276
rect 38332 15426 38388 15484
rect 38332 15374 38334 15426
rect 38386 15374 38388 15426
rect 38332 15362 38388 15374
rect 38444 15986 38612 15988
rect 38444 15934 38558 15986
rect 38610 15934 38612 15986
rect 38444 15932 38612 15934
rect 38220 15262 38222 15314
rect 38274 15262 38276 15314
rect 38220 15250 38276 15262
rect 38444 15148 38500 15932
rect 38556 15922 38612 15932
rect 38668 17220 38724 17230
rect 38108 15092 38276 15148
rect 37996 14702 37998 14754
rect 38050 14702 38052 14754
rect 37996 14690 38052 14702
rect 38108 14980 38164 14990
rect 37884 14476 38052 14532
rect 37660 14420 37716 14430
rect 37716 14364 37828 14420
rect 37660 14326 37716 14364
rect 37548 13524 37604 13534
rect 37548 13430 37604 13468
rect 37772 13524 37828 14364
rect 37884 14308 37940 14318
rect 37884 14214 37940 14252
rect 37548 13188 37604 13198
rect 37548 13074 37604 13132
rect 37548 13022 37550 13074
rect 37602 13022 37604 13074
rect 37548 13010 37604 13022
rect 37660 12964 37716 12974
rect 37772 12964 37828 13468
rect 37884 12964 37940 12974
rect 37772 12962 37940 12964
rect 37772 12910 37886 12962
rect 37938 12910 37940 12962
rect 37772 12908 37940 12910
rect 37324 12292 37380 12302
rect 37324 12198 37380 12236
rect 37548 12178 37604 12190
rect 37548 12126 37550 12178
rect 37602 12126 37604 12178
rect 37548 11394 37604 12126
rect 37660 11508 37716 12908
rect 37884 12898 37940 12908
rect 37996 12740 38052 14476
rect 37772 12684 38052 12740
rect 37772 12402 37828 12684
rect 37772 12350 37774 12402
rect 37826 12350 37828 12402
rect 37772 11732 37828 12350
rect 37772 11666 37828 11676
rect 37884 12178 37940 12190
rect 37884 12126 37886 12178
rect 37938 12126 37940 12178
rect 37660 11452 37828 11508
rect 37548 11342 37550 11394
rect 37602 11342 37604 11394
rect 37548 11330 37604 11342
rect 37212 10782 37214 10834
rect 37266 10782 37268 10834
rect 37212 10770 37268 10782
rect 37100 10658 37156 10668
rect 37660 10724 37716 10734
rect 37660 10610 37716 10668
rect 37660 10558 37662 10610
rect 37714 10558 37716 10610
rect 37660 10546 37716 10558
rect 35868 9102 35870 9154
rect 35922 9102 35924 9154
rect 35868 9090 35924 9102
rect 36204 9324 36372 9380
rect 36540 10332 36820 10388
rect 36204 8932 36260 9324
rect 36204 8866 36260 8876
rect 36316 9042 36372 9054
rect 36316 8990 36318 9042
rect 36370 8990 36372 9042
rect 35308 8764 35588 8820
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35532 8484 35588 8764
rect 35084 7646 35086 7698
rect 35138 7646 35140 7698
rect 35084 7634 35140 7646
rect 35420 8428 35588 8484
rect 35420 7476 35476 8428
rect 35644 8372 35700 8382
rect 35644 8258 35700 8316
rect 35644 8206 35646 8258
rect 35698 8206 35700 8258
rect 35644 8194 35700 8206
rect 36204 8372 36260 8382
rect 35868 8034 35924 8046
rect 35868 7982 35870 8034
rect 35922 7982 35924 8034
rect 34804 7420 34916 7476
rect 35084 7420 35476 7476
rect 35532 7586 35588 7598
rect 35532 7534 35534 7586
rect 35586 7534 35588 7586
rect 34748 6580 34804 7420
rect 34636 6578 34804 6580
rect 34636 6526 34750 6578
rect 34802 6526 34804 6578
rect 34636 6524 34804 6526
rect 34524 6468 34580 6478
rect 34524 6374 34580 6412
rect 34132 6076 34356 6132
rect 34076 5906 34132 6076
rect 34636 6020 34692 6524
rect 34748 6514 34804 6524
rect 34972 7364 35028 7374
rect 34076 5854 34078 5906
rect 34130 5854 34132 5906
rect 34076 5842 34132 5854
rect 34300 5964 34916 6020
rect 33852 5628 34244 5684
rect 33516 5516 33684 5572
rect 33292 5236 33348 5246
rect 33292 5142 33348 5180
rect 33180 4946 33236 4956
rect 33180 4788 33236 4798
rect 33180 4562 33236 4732
rect 33180 4510 33182 4562
rect 33234 4510 33236 4562
rect 33180 4498 33236 4510
rect 33628 4226 33684 5516
rect 33740 5124 33796 5134
rect 33740 5030 33796 5068
rect 34188 4562 34244 5628
rect 34300 5234 34356 5964
rect 34300 5182 34302 5234
rect 34354 5182 34356 5234
rect 34300 5170 34356 5182
rect 34860 5236 34916 5964
rect 34972 5906 35028 7308
rect 35084 6916 35140 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 6916 35252 6926
rect 35084 6860 35196 6916
rect 35196 6690 35252 6860
rect 35532 6914 35588 7534
rect 35644 7364 35700 7374
rect 35644 7270 35700 7308
rect 35756 7252 35812 7262
rect 35868 7252 35924 7982
rect 36092 7362 36148 7374
rect 36092 7310 36094 7362
rect 36146 7310 36148 7362
rect 36092 7252 36148 7310
rect 35756 7250 36148 7252
rect 35756 7198 35758 7250
rect 35810 7198 36148 7250
rect 35756 7196 36148 7198
rect 35756 7186 35812 7196
rect 35532 6862 35534 6914
rect 35586 6862 35588 6914
rect 35532 6850 35588 6862
rect 35196 6638 35198 6690
rect 35250 6638 35252 6690
rect 35196 6626 35252 6638
rect 35644 6466 35700 6478
rect 35644 6414 35646 6466
rect 35698 6414 35700 6466
rect 35644 6244 35700 6414
rect 35700 6188 36036 6244
rect 35644 6178 35700 6188
rect 35980 6130 36036 6188
rect 35980 6078 35982 6130
rect 36034 6078 36036 6130
rect 35980 6066 36036 6078
rect 35196 6020 35252 6030
rect 35196 5926 35252 5964
rect 34972 5854 34974 5906
rect 35026 5854 35028 5906
rect 34972 5842 35028 5854
rect 36092 5684 36148 7196
rect 36204 6802 36260 8316
rect 36316 8148 36372 8990
rect 36316 8054 36372 8092
rect 36540 7588 36596 10332
rect 37772 10052 37828 11452
rect 37884 11172 37940 12126
rect 37996 11396 38052 11406
rect 37996 11302 38052 11340
rect 37884 11106 37940 11116
rect 37772 9996 37940 10052
rect 37100 9940 37156 9950
rect 37100 9846 37156 9884
rect 37436 9826 37492 9838
rect 37436 9774 37438 9826
rect 37490 9774 37492 9826
rect 36988 9154 37044 9166
rect 36988 9102 36990 9154
rect 37042 9102 37044 9154
rect 36764 9042 36820 9054
rect 36764 8990 36766 9042
rect 36818 8990 36820 9042
rect 36652 7700 36708 7710
rect 36652 7606 36708 7644
rect 36540 7522 36596 7532
rect 36204 6750 36206 6802
rect 36258 6750 36260 6802
rect 36204 6738 36260 6750
rect 36316 7252 36372 7262
rect 36764 7252 36820 8990
rect 36988 8372 37044 9102
rect 36988 8306 37044 8316
rect 37100 9156 37156 9166
rect 37100 8258 37156 9100
rect 37436 8370 37492 9774
rect 37436 8318 37438 8370
rect 37490 8318 37492 8370
rect 37436 8306 37492 8318
rect 37884 8372 37940 9996
rect 37996 9828 38052 9838
rect 37996 9734 38052 9772
rect 38108 9156 38164 14924
rect 38220 12964 38276 15092
rect 38220 12898 38276 12908
rect 38332 15092 38500 15148
rect 38556 15204 38612 15214
rect 38332 14084 38388 15092
rect 38332 12852 38388 14028
rect 38444 14420 38500 14430
rect 38444 13746 38500 14364
rect 38444 13694 38446 13746
rect 38498 13694 38500 13746
rect 38444 13076 38500 13694
rect 38444 13010 38500 13020
rect 38556 13524 38612 15148
rect 38668 15202 38724 17164
rect 39004 17108 39060 17502
rect 38892 17052 39060 17108
rect 39116 17444 39172 17454
rect 38668 15150 38670 15202
rect 38722 15150 38724 15202
rect 38668 15138 38724 15150
rect 38780 16770 38836 16782
rect 38780 16718 38782 16770
rect 38834 16718 38836 16770
rect 38780 15148 38836 16718
rect 38892 16772 38948 17052
rect 39116 16996 39172 17388
rect 39116 16882 39172 16940
rect 39116 16830 39118 16882
rect 39170 16830 39172 16882
rect 39116 16818 39172 16830
rect 38892 15652 38948 16716
rect 38892 15586 38948 15596
rect 39228 15316 39284 17612
rect 39340 17602 39396 17612
rect 39564 17108 39620 18284
rect 39676 20578 39844 20580
rect 39676 20526 39790 20578
rect 39842 20526 39844 20578
rect 39676 20524 39844 20526
rect 39676 18116 39732 20524
rect 39788 20514 39844 20524
rect 40012 19684 40068 19694
rect 39788 18452 39844 18462
rect 39788 18358 39844 18396
rect 39676 18050 39732 18060
rect 39900 17668 39956 17678
rect 39676 17444 39732 17454
rect 39676 17350 39732 17388
rect 39676 17108 39732 17118
rect 39564 17106 39732 17108
rect 39564 17054 39678 17106
rect 39730 17054 39732 17106
rect 39564 17052 39732 17054
rect 39676 17042 39732 17052
rect 39788 17108 39844 17118
rect 39564 16882 39620 16894
rect 39564 16830 39566 16882
rect 39618 16830 39620 16882
rect 39564 16212 39620 16830
rect 39564 16098 39620 16156
rect 39564 16046 39566 16098
rect 39618 16046 39620 16098
rect 39564 16034 39620 16046
rect 39004 15314 39284 15316
rect 39004 15262 39230 15314
rect 39282 15262 39284 15314
rect 39004 15260 39284 15262
rect 38780 15092 38948 15148
rect 38668 14756 38724 14766
rect 38668 14530 38724 14700
rect 38668 14478 38670 14530
rect 38722 14478 38724 14530
rect 38668 13748 38724 14478
rect 38892 14418 38948 15092
rect 38892 14366 38894 14418
rect 38946 14366 38948 14418
rect 38892 14354 38948 14366
rect 38668 13682 38724 13692
rect 38892 13634 38948 13646
rect 38892 13582 38894 13634
rect 38946 13582 38948 13634
rect 38668 13524 38724 13534
rect 38556 13522 38724 13524
rect 38556 13470 38670 13522
rect 38722 13470 38724 13522
rect 38556 13468 38724 13470
rect 38556 12964 38612 13468
rect 38668 13458 38724 13468
rect 38892 13524 38948 13582
rect 38556 12908 38724 12964
rect 38444 12852 38500 12862
rect 38332 12850 38500 12852
rect 38332 12798 38446 12850
rect 38498 12798 38500 12850
rect 38332 12796 38500 12798
rect 38444 12786 38500 12796
rect 38220 12740 38276 12750
rect 38220 12404 38276 12684
rect 38556 12740 38612 12750
rect 38556 12646 38612 12684
rect 38220 12338 38276 12348
rect 38444 12404 38500 12414
rect 38668 12404 38724 12908
rect 38444 12402 38724 12404
rect 38444 12350 38446 12402
rect 38498 12350 38724 12402
rect 38444 12348 38724 12350
rect 38892 12404 38948 13468
rect 39004 12964 39060 15260
rect 39228 15250 39284 15260
rect 39340 15874 39396 15886
rect 39340 15822 39342 15874
rect 39394 15822 39396 15874
rect 39340 14980 39396 15822
rect 39340 14914 39396 14924
rect 39788 15538 39844 17052
rect 39900 17106 39956 17612
rect 39900 17054 39902 17106
rect 39954 17054 39956 17106
rect 39900 17042 39956 17054
rect 39788 15486 39790 15538
rect 39842 15486 39844 15538
rect 39788 14868 39844 15486
rect 39788 14802 39844 14812
rect 39900 16098 39956 16110
rect 39900 16046 39902 16098
rect 39954 16046 39956 16098
rect 39900 14756 39956 16046
rect 39900 14690 39956 14700
rect 40012 14308 40068 19628
rect 40124 17442 40180 17454
rect 40124 17390 40126 17442
rect 40178 17390 40180 17442
rect 40124 16772 40180 17390
rect 40124 16706 40180 16716
rect 40348 16772 40404 23548
rect 40796 22708 40852 23886
rect 41244 23714 41300 25228
rect 41244 23662 41246 23714
rect 41298 23662 41300 23714
rect 41244 23650 41300 23662
rect 41804 24834 41860 24846
rect 41804 24782 41806 24834
rect 41858 24782 41860 24834
rect 41804 23716 41860 24782
rect 41916 24724 41972 26460
rect 42140 26450 42196 26460
rect 42364 25844 42420 28364
rect 42812 28326 42868 28364
rect 43260 27636 43316 27646
rect 43260 27298 43316 27580
rect 43260 27246 43262 27298
rect 43314 27246 43316 27298
rect 43260 27234 43316 27246
rect 43372 27076 43428 28478
rect 43484 28532 43540 28542
rect 43596 28532 43652 28588
rect 43932 28578 43988 28588
rect 43484 28530 43652 28532
rect 43484 28478 43486 28530
rect 43538 28478 43652 28530
rect 43484 28476 43652 28478
rect 44492 28532 44548 29486
rect 45276 29204 45332 29214
rect 45276 29110 45332 29148
rect 45052 28644 45108 28654
rect 45052 28642 45220 28644
rect 45052 28590 45054 28642
rect 45106 28590 45220 28642
rect 45052 28588 45220 28590
rect 45052 28578 45108 28588
rect 43484 27188 43540 28476
rect 44492 28082 44548 28476
rect 44492 28030 44494 28082
rect 44546 28030 44548 28082
rect 44492 28018 44548 28030
rect 45164 28420 45220 28588
rect 45164 27748 45220 28364
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 46396 27970 46452 27982
rect 46396 27918 46398 27970
rect 46450 27918 46452 27970
rect 45388 27748 45444 27758
rect 45836 27748 45892 27758
rect 45164 27746 45444 27748
rect 45164 27694 45390 27746
rect 45442 27694 45444 27746
rect 45164 27692 45444 27694
rect 45052 27636 45108 27646
rect 45052 27542 45108 27580
rect 43596 27188 43652 27198
rect 43484 27132 43596 27188
rect 43596 27122 43652 27132
rect 43372 27020 43540 27076
rect 43484 26962 43540 27020
rect 43484 26910 43486 26962
rect 43538 26910 43540 26962
rect 43484 26898 43540 26910
rect 43596 26964 43652 26974
rect 43372 26850 43428 26862
rect 43372 26798 43374 26850
rect 43426 26798 43428 26850
rect 43372 26740 43428 26798
rect 43260 26684 43428 26740
rect 43036 26404 43092 26414
rect 42140 25788 42420 25844
rect 42588 26402 43092 26404
rect 42588 26350 43038 26402
rect 43090 26350 43092 26402
rect 42588 26348 43092 26350
rect 42140 24948 42196 25788
rect 42364 25620 42420 25630
rect 42364 25506 42420 25564
rect 42588 25618 42644 26348
rect 43036 26338 43092 26348
rect 43148 26402 43204 26414
rect 43148 26350 43150 26402
rect 43202 26350 43204 26402
rect 43148 26292 43204 26350
rect 42700 26178 42756 26190
rect 42700 26126 42702 26178
rect 42754 26126 42756 26178
rect 42700 25956 42756 26126
rect 43148 25956 43204 26236
rect 42700 25900 43204 25956
rect 42588 25566 42590 25618
rect 42642 25566 42644 25618
rect 42588 25554 42644 25566
rect 42364 25454 42366 25506
rect 42418 25454 42420 25506
rect 42364 25396 42420 25454
rect 42364 25330 42420 25340
rect 42700 25506 42756 25518
rect 42700 25454 42702 25506
rect 42754 25454 42756 25506
rect 42140 24946 42532 24948
rect 42140 24894 42142 24946
rect 42194 24894 42532 24946
rect 42140 24892 42532 24894
rect 42140 24882 42196 24892
rect 41916 24668 42308 24724
rect 42028 23716 42084 23726
rect 41804 23660 42028 23716
rect 42028 23622 42084 23660
rect 41020 23268 41076 23278
rect 41020 23174 41076 23212
rect 41804 23268 41860 23278
rect 41804 23174 41860 23212
rect 40908 23156 40964 23166
rect 40908 23062 40964 23100
rect 42140 23044 42196 23054
rect 42140 22950 42196 22988
rect 40796 22642 40852 22652
rect 41020 22820 41076 22830
rect 41020 21698 41076 22764
rect 41916 22820 41972 22830
rect 41972 22764 42084 22820
rect 41916 22754 41972 22764
rect 41356 22370 41412 22382
rect 41580 22372 41636 22382
rect 41356 22318 41358 22370
rect 41410 22318 41412 22370
rect 41020 21646 41022 21698
rect 41074 21646 41076 21698
rect 41020 21634 41076 21646
rect 41132 22148 41188 22158
rect 40460 21476 40516 21486
rect 40460 20690 40516 21420
rect 40460 20638 40462 20690
rect 40514 20638 40516 20690
rect 40460 20626 40516 20638
rect 40572 20692 40628 20702
rect 40572 20598 40628 20636
rect 41132 20468 41188 22092
rect 41244 21476 41300 21486
rect 41244 21382 41300 21420
rect 41356 20804 41412 22318
rect 41468 22370 41636 22372
rect 41468 22318 41582 22370
rect 41634 22318 41636 22370
rect 41468 22316 41636 22318
rect 41468 21476 41524 22316
rect 41580 22306 41636 22316
rect 42028 22370 42084 22764
rect 42028 22318 42030 22370
rect 42082 22318 42084 22370
rect 42028 22306 42084 22318
rect 41468 21410 41524 21420
rect 41804 22258 41860 22270
rect 41804 22206 41806 22258
rect 41858 22206 41860 22258
rect 41580 21364 41636 21374
rect 41804 21364 41860 22206
rect 42140 22260 42196 22270
rect 42252 22260 42308 24668
rect 42476 24050 42532 24892
rect 42476 23998 42478 24050
rect 42530 23998 42532 24050
rect 42476 23986 42532 23998
rect 42588 24836 42644 24846
rect 42700 24836 42756 25454
rect 42644 24780 42756 24836
rect 42588 23714 42644 24780
rect 42588 23662 42590 23714
rect 42642 23662 42644 23714
rect 42364 23266 42420 23278
rect 42364 23214 42366 23266
rect 42418 23214 42420 23266
rect 42364 22820 42420 23214
rect 42364 22754 42420 22764
rect 42140 22258 42308 22260
rect 42140 22206 42142 22258
rect 42194 22206 42308 22258
rect 42140 22204 42308 22206
rect 42140 21812 42196 22204
rect 42140 21746 42196 21756
rect 42252 21698 42308 21710
rect 42252 21646 42254 21698
rect 42306 21646 42308 21698
rect 42140 21586 42196 21598
rect 42140 21534 42142 21586
rect 42194 21534 42196 21586
rect 41916 21364 41972 21374
rect 41580 21362 41748 21364
rect 41580 21310 41582 21362
rect 41634 21310 41748 21362
rect 41580 21308 41748 21310
rect 41804 21308 41916 21364
rect 41580 21298 41636 21308
rect 41580 20804 41636 20814
rect 41356 20802 41636 20804
rect 41356 20750 41582 20802
rect 41634 20750 41636 20802
rect 41356 20748 41636 20750
rect 41580 20692 41636 20748
rect 41580 20626 41636 20636
rect 41692 20690 41748 21308
rect 41916 21298 41972 21308
rect 41692 20638 41694 20690
rect 41746 20638 41748 20690
rect 41692 20626 41748 20638
rect 42140 20692 42196 21534
rect 42140 20626 42196 20636
rect 42252 21476 42308 21646
rect 41692 20468 41748 20478
rect 41132 20412 41636 20468
rect 41580 20018 41636 20412
rect 41580 19966 41582 20018
rect 41634 19966 41636 20018
rect 41580 19458 41636 19966
rect 41580 19406 41582 19458
rect 41634 19406 41636 19458
rect 41580 19394 41636 19406
rect 41692 19236 41748 20412
rect 41916 20018 41972 20030
rect 41916 19966 41918 20018
rect 41970 19966 41972 20018
rect 41804 19908 41860 19918
rect 41804 19814 41860 19852
rect 41916 19684 41972 19966
rect 41580 19180 41748 19236
rect 41804 19628 41972 19684
rect 42140 20018 42196 20030
rect 42140 19966 42142 20018
rect 42194 19966 42196 20018
rect 41804 19236 41860 19628
rect 42140 19572 42196 19966
rect 41916 19516 42196 19572
rect 41916 19458 41972 19516
rect 41916 19406 41918 19458
rect 41970 19406 41972 19458
rect 41916 19394 41972 19406
rect 41804 19180 41972 19236
rect 41244 18562 41300 18574
rect 41244 18510 41246 18562
rect 41298 18510 41300 18562
rect 41020 18450 41076 18462
rect 41020 18398 41022 18450
rect 41074 18398 41076 18450
rect 41020 17780 41076 18398
rect 41020 17714 41076 17724
rect 40348 16706 40404 16716
rect 40908 17666 40964 17678
rect 40908 17614 40910 17666
rect 40962 17614 40964 17666
rect 40908 16660 40964 17614
rect 41132 17556 41188 17566
rect 41132 17462 41188 17500
rect 41244 17444 41300 18510
rect 41244 17378 41300 17388
rect 41468 16994 41524 17006
rect 41468 16942 41470 16994
rect 41522 16942 41524 16994
rect 41356 16882 41412 16894
rect 41356 16830 41358 16882
rect 41410 16830 41412 16882
rect 41356 16772 41412 16830
rect 41468 16884 41524 16942
rect 41468 16818 41524 16828
rect 41356 16706 41412 16716
rect 40908 16594 40964 16604
rect 41580 16548 41636 19180
rect 41804 19010 41860 19022
rect 41804 18958 41806 19010
rect 41858 18958 41860 19010
rect 41804 18452 41860 18958
rect 41804 18226 41860 18396
rect 41916 18340 41972 19180
rect 42140 19012 42196 19022
rect 42140 18450 42196 18956
rect 42140 18398 42142 18450
rect 42194 18398 42196 18450
rect 42140 18386 42196 18398
rect 41916 18274 41972 18284
rect 41804 18174 41806 18226
rect 41858 18174 41860 18226
rect 41692 17666 41748 17678
rect 41692 17614 41694 17666
rect 41746 17614 41748 17666
rect 41692 17444 41748 17614
rect 41804 17556 41860 18174
rect 41804 17490 41860 17500
rect 41692 17378 41748 17388
rect 42028 17444 42084 17454
rect 42028 17350 42084 17388
rect 41916 17332 41972 17342
rect 41356 16492 41636 16548
rect 41804 16772 41860 16782
rect 40348 16324 40404 16334
rect 40236 15202 40292 15214
rect 40236 15150 40238 15202
rect 40290 15150 40292 15202
rect 40236 15148 40292 15150
rect 40124 15092 40292 15148
rect 40348 15148 40404 16268
rect 41244 15204 41300 15242
rect 40348 15092 40516 15148
rect 41244 15138 41300 15148
rect 40124 14420 40180 15092
rect 40236 14980 40292 14990
rect 40236 14530 40292 14924
rect 40236 14478 40238 14530
rect 40290 14478 40292 14530
rect 40236 14466 40292 14478
rect 40124 14354 40180 14364
rect 39788 14252 40068 14308
rect 39004 12962 39396 12964
rect 39004 12910 39006 12962
rect 39058 12910 39396 12962
rect 39004 12908 39396 12910
rect 39004 12898 39060 12908
rect 38892 12348 39060 12404
rect 38444 12338 38500 12348
rect 38892 12178 38948 12190
rect 38892 12126 38894 12178
rect 38946 12126 38948 12178
rect 38780 11732 38836 11742
rect 38444 11508 38500 11518
rect 38444 11414 38500 11452
rect 38780 11282 38836 11676
rect 38780 11230 38782 11282
rect 38834 11230 38836 11282
rect 38780 11218 38836 11230
rect 38892 11506 38948 12126
rect 38892 11454 38894 11506
rect 38946 11454 38948 11506
rect 38332 11170 38388 11182
rect 38332 11118 38334 11170
rect 38386 11118 38388 11170
rect 38108 9090 38164 9100
rect 38220 10722 38276 10734
rect 38220 10670 38222 10722
rect 38274 10670 38276 10722
rect 38220 10500 38276 10670
rect 38332 10724 38388 11118
rect 38332 10658 38388 10668
rect 38556 11172 38612 11182
rect 38556 10500 38612 11116
rect 38220 10444 38612 10500
rect 38220 8930 38276 10444
rect 38220 8878 38222 8930
rect 38274 8878 38276 8930
rect 38220 8866 38276 8878
rect 38556 9940 38612 9950
rect 38556 8428 38612 9884
rect 38892 9940 38948 11454
rect 38892 9874 38948 9884
rect 39004 11060 39060 12348
rect 39340 12402 39396 12908
rect 39676 12962 39732 12974
rect 39676 12910 39678 12962
rect 39730 12910 39732 12962
rect 39340 12350 39342 12402
rect 39394 12350 39396 12402
rect 39340 12338 39396 12350
rect 39452 12740 39508 12750
rect 39452 12402 39508 12684
rect 39452 12350 39454 12402
rect 39506 12350 39508 12402
rect 39452 12338 39508 12350
rect 39564 12180 39620 12190
rect 39564 12086 39620 12124
rect 39676 11618 39732 12910
rect 39676 11566 39678 11618
rect 39730 11566 39732 11618
rect 39676 11554 39732 11566
rect 39340 11170 39396 11182
rect 39340 11118 39342 11170
rect 39394 11118 39396 11170
rect 39340 11060 39396 11118
rect 39004 11004 39396 11060
rect 38780 9156 38836 9166
rect 38780 9062 38836 9100
rect 37996 8372 38052 8382
rect 38556 8372 38836 8428
rect 37940 8370 38052 8372
rect 37940 8318 37998 8370
rect 38050 8318 38052 8370
rect 37940 8316 38052 8318
rect 37884 8278 37940 8316
rect 37996 8306 38052 8316
rect 37100 8206 37102 8258
rect 37154 8206 37156 8258
rect 37100 8194 37156 8206
rect 37212 8148 37268 8158
rect 37212 7588 37268 8092
rect 37548 8146 37604 8158
rect 37548 8094 37550 8146
rect 37602 8094 37604 8146
rect 37548 7700 37604 8094
rect 38444 8148 38500 8158
rect 38444 8054 38500 8092
rect 36316 7250 36820 7252
rect 36316 7198 36318 7250
rect 36370 7198 36820 7250
rect 36316 7196 36820 7198
rect 36876 7532 37380 7588
rect 36316 6244 36372 7196
rect 36316 6178 36372 6188
rect 36540 6914 36596 6926
rect 36540 6862 36542 6914
rect 36594 6862 36596 6914
rect 36540 6580 36596 6862
rect 36540 6130 36596 6524
rect 36540 6078 36542 6130
rect 36594 6078 36596 6130
rect 36540 6066 36596 6078
rect 36092 5618 36148 5628
rect 36876 5794 36932 7532
rect 37324 7474 37380 7532
rect 37324 7422 37326 7474
rect 37378 7422 37380 7474
rect 37324 7410 37380 7422
rect 37100 7364 37156 7374
rect 37100 6802 37156 7308
rect 37548 7252 37604 7644
rect 38444 7588 38500 7598
rect 37884 7586 38500 7588
rect 37884 7534 38446 7586
rect 38498 7534 38500 7586
rect 37884 7532 38500 7534
rect 37884 7474 37940 7532
rect 38444 7522 38500 7532
rect 37884 7422 37886 7474
rect 37938 7422 37940 7474
rect 37884 7410 37940 7422
rect 38668 7476 38724 7486
rect 37996 7364 38052 7374
rect 37996 7270 38052 7308
rect 37548 7186 37604 7196
rect 38332 7252 38388 7262
rect 38332 7158 38388 7196
rect 37100 6750 37102 6802
rect 37154 6750 37156 6802
rect 37100 6738 37156 6750
rect 37324 6690 37380 6702
rect 37324 6638 37326 6690
rect 37378 6638 37380 6690
rect 37324 6244 37380 6638
rect 37996 6692 38052 6702
rect 38668 6692 38724 7420
rect 37996 6598 38052 6636
rect 38444 6636 38724 6692
rect 38444 6580 38500 6636
rect 38444 6486 38500 6524
rect 37324 6130 37380 6188
rect 37324 6078 37326 6130
rect 37378 6078 37380 6130
rect 37324 6066 37380 6078
rect 36876 5742 36878 5794
rect 36930 5742 36932 5794
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35420 5348 35476 5358
rect 35084 5236 35140 5246
rect 34860 5234 35140 5236
rect 34860 5182 35086 5234
rect 35138 5182 35140 5234
rect 34860 5180 35140 5182
rect 35084 5170 35140 5180
rect 35420 5234 35476 5292
rect 35420 5182 35422 5234
rect 35474 5182 35476 5234
rect 35420 5170 35476 5182
rect 34188 4510 34190 4562
rect 34242 4510 34244 4562
rect 34188 4498 34244 4510
rect 34524 4564 34580 4574
rect 34524 4470 34580 4508
rect 33628 4174 33630 4226
rect 33682 4174 33684 4226
rect 33628 4162 33684 4174
rect 35196 3948 35460 3958
rect 33180 3892 33236 3902
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 33180 3668 33236 3836
rect 33628 3668 33684 3678
rect 33180 3666 33684 3668
rect 33180 3614 33182 3666
rect 33234 3614 33630 3666
rect 33682 3614 33684 3666
rect 33180 3612 33684 3614
rect 33180 3602 33236 3612
rect 33628 3602 33684 3612
rect 34076 3668 34132 3678
rect 34076 3574 34132 3612
rect 32732 3332 32788 3342
rect 32732 3238 32788 3276
rect 36876 2660 36932 5742
rect 38780 3108 38836 8372
rect 38892 5684 38948 5694
rect 38892 5234 38948 5628
rect 38892 5182 38894 5234
rect 38946 5182 38948 5234
rect 38892 5170 38948 5182
rect 38780 3042 38836 3052
rect 36876 2594 36932 2604
rect 32508 2370 32564 2380
rect 26908 1586 26964 1596
rect 39004 1540 39060 11004
rect 39788 10276 39844 14252
rect 40012 14084 40068 14094
rect 39900 13748 39956 13758
rect 39900 13654 39956 13692
rect 40012 13746 40068 14028
rect 40012 13694 40014 13746
rect 40066 13694 40068 13746
rect 40012 13682 40068 13694
rect 40460 12964 40516 15092
rect 41020 14868 41076 14878
rect 41020 14530 41076 14812
rect 41020 14478 41022 14530
rect 41074 14478 41076 14530
rect 41020 14466 41076 14478
rect 40796 14418 40852 14430
rect 40796 14366 40798 14418
rect 40850 14366 40852 14418
rect 40012 12852 40068 12862
rect 39900 12404 39956 12414
rect 39900 11506 39956 12348
rect 40012 12290 40068 12796
rect 40124 12740 40180 12750
rect 40124 12402 40180 12684
rect 40124 12350 40126 12402
rect 40178 12350 40180 12402
rect 40124 12338 40180 12350
rect 40012 12238 40014 12290
rect 40066 12238 40068 12290
rect 40012 12226 40068 12238
rect 39900 11454 39902 11506
rect 39954 11454 39956 11506
rect 39900 11442 39956 11454
rect 40124 11954 40180 11966
rect 40124 11902 40126 11954
rect 40178 11902 40180 11954
rect 39452 10220 39844 10276
rect 39900 10836 39956 10846
rect 39340 9716 39396 9726
rect 39340 9622 39396 9660
rect 39116 9268 39172 9278
rect 39452 9268 39508 10220
rect 39564 10052 39620 10062
rect 39564 9826 39620 9996
rect 39564 9774 39566 9826
rect 39618 9774 39620 9826
rect 39564 9762 39620 9774
rect 39900 9828 39956 10780
rect 40124 10164 40180 11902
rect 40236 11618 40292 11630
rect 40236 11566 40238 11618
rect 40290 11566 40292 11618
rect 40236 11506 40292 11566
rect 40460 11618 40516 12908
rect 40460 11566 40462 11618
rect 40514 11566 40516 11618
rect 40460 11554 40516 11566
rect 40684 13076 40740 13086
rect 40684 12962 40740 13020
rect 40684 12910 40686 12962
rect 40738 12910 40740 12962
rect 40684 12180 40740 12910
rect 40796 12628 40852 14366
rect 40908 13636 40964 13646
rect 40908 13074 40964 13580
rect 41020 13634 41076 13646
rect 41020 13582 41022 13634
rect 41074 13582 41076 13634
rect 41020 13524 41076 13582
rect 41020 13458 41076 13468
rect 40908 13022 40910 13074
rect 40962 13022 40964 13074
rect 40908 13010 40964 13022
rect 40796 12562 40852 12572
rect 41244 12516 41300 12526
rect 41244 12290 41300 12460
rect 41244 12238 41246 12290
rect 41298 12238 41300 12290
rect 41244 12226 41300 12238
rect 40236 11454 40238 11506
rect 40290 11454 40292 11506
rect 40236 11442 40292 11454
rect 40684 11170 40740 12124
rect 41244 11618 41300 11630
rect 41244 11566 41246 11618
rect 41298 11566 41300 11618
rect 41244 11506 41300 11566
rect 41244 11454 41246 11506
rect 41298 11454 41300 11506
rect 41244 11442 41300 11454
rect 40684 11118 40686 11170
rect 40738 11118 40740 11170
rect 40124 10108 40404 10164
rect 40348 10052 40404 10108
rect 40348 9996 40516 10052
rect 39900 9826 40292 9828
rect 39900 9774 39902 9826
rect 39954 9774 40292 9826
rect 39900 9772 40292 9774
rect 39900 9762 39956 9772
rect 39564 9604 39620 9614
rect 39564 9602 39956 9604
rect 39564 9550 39566 9602
rect 39618 9550 39956 9602
rect 39564 9548 39956 9550
rect 39564 9538 39620 9548
rect 39564 9268 39620 9278
rect 39116 9266 39620 9268
rect 39116 9214 39118 9266
rect 39170 9214 39566 9266
rect 39618 9214 39620 9266
rect 39116 9212 39620 9214
rect 39116 7476 39172 9212
rect 39564 9202 39620 9212
rect 39116 7410 39172 7420
rect 39340 9044 39396 9054
rect 39340 7474 39396 8988
rect 39900 8260 39956 9548
rect 40236 9266 40292 9772
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 40236 9202 40292 9214
rect 40348 9826 40404 9838
rect 40348 9774 40350 9826
rect 40402 9774 40404 9826
rect 39900 8194 39956 8204
rect 40348 8258 40404 9774
rect 40348 8206 40350 8258
rect 40402 8206 40404 8258
rect 39340 7422 39342 7474
rect 39394 7422 39396 7474
rect 39116 6468 39172 6478
rect 39340 6468 39396 7422
rect 39564 7362 39620 7374
rect 39564 7310 39566 7362
rect 39618 7310 39620 7362
rect 39564 6580 39620 7310
rect 39676 7364 39732 7374
rect 40124 7364 40180 7374
rect 39676 7362 40180 7364
rect 39676 7310 39678 7362
rect 39730 7310 40126 7362
rect 40178 7310 40180 7362
rect 39676 7308 40180 7310
rect 39676 7298 39732 7308
rect 40124 6804 40180 7308
rect 40236 6804 40292 6814
rect 40124 6748 40236 6804
rect 40236 6738 40292 6748
rect 39564 6524 40292 6580
rect 39116 6466 39396 6468
rect 39116 6414 39118 6466
rect 39170 6414 39396 6466
rect 39116 6412 39396 6414
rect 39116 3220 39172 6412
rect 40236 6018 40292 6524
rect 40348 6468 40404 8206
rect 40460 6804 40516 9996
rect 40572 9716 40628 9726
rect 40572 8932 40628 9660
rect 40684 9156 40740 11118
rect 41356 10836 41412 16492
rect 41468 16098 41524 16110
rect 41468 16046 41470 16098
rect 41522 16046 41524 16098
rect 41468 15316 41524 16046
rect 41468 15250 41524 15260
rect 41804 13858 41860 16716
rect 41916 16660 41972 17276
rect 41916 16594 41972 16604
rect 42140 16884 42196 16894
rect 42028 16548 42084 16558
rect 42028 16436 42084 16492
rect 41916 16380 42084 16436
rect 41916 14530 41972 16380
rect 42140 16210 42196 16828
rect 42140 16158 42142 16210
rect 42194 16158 42196 16210
rect 42140 16146 42196 16158
rect 42252 15988 42308 21420
rect 42476 21364 42532 21374
rect 42476 20802 42532 21308
rect 42476 20750 42478 20802
rect 42530 20750 42532 20802
rect 42476 20738 42532 20750
rect 42476 20580 42532 20590
rect 42364 20578 42532 20580
rect 42364 20526 42478 20578
rect 42530 20526 42532 20578
rect 42364 20524 42532 20526
rect 42364 16772 42420 20524
rect 42476 20514 42532 20524
rect 42588 20356 42644 23662
rect 42700 23716 42756 23726
rect 42700 23154 42756 23660
rect 42812 23268 42868 25900
rect 43260 25844 43316 26684
rect 43372 26516 43428 26526
rect 43596 26516 43652 26908
rect 43372 26514 43652 26516
rect 43372 26462 43374 26514
rect 43426 26462 43652 26514
rect 43372 26460 43652 26462
rect 43372 26450 43428 26460
rect 43708 26292 43764 26302
rect 43708 26198 43764 26236
rect 42812 23202 42868 23212
rect 42924 25788 43316 25844
rect 42700 23102 42702 23154
rect 42754 23102 42756 23154
rect 42700 21588 42756 23102
rect 42812 21924 42868 21934
rect 42812 21810 42868 21868
rect 42812 21758 42814 21810
rect 42866 21758 42868 21810
rect 42812 21746 42868 21758
rect 42812 21588 42868 21598
rect 42700 21532 42812 21588
rect 42812 20468 42868 21532
rect 42812 20402 42868 20412
rect 42476 20300 42644 20356
rect 42476 17220 42532 20300
rect 42924 19348 42980 25788
rect 43484 25620 43540 25630
rect 43036 25618 43540 25620
rect 43036 25566 43486 25618
rect 43538 25566 43540 25618
rect 43036 25564 43540 25566
rect 43036 25506 43092 25564
rect 43484 25554 43540 25564
rect 43036 25454 43038 25506
rect 43090 25454 43092 25506
rect 43036 25442 43092 25454
rect 45164 25508 45220 25518
rect 43372 25396 43428 25406
rect 43372 25302 43428 25340
rect 43596 25282 43652 25294
rect 43596 25230 43598 25282
rect 43650 25230 43652 25282
rect 43372 24836 43428 24846
rect 43372 24742 43428 24780
rect 43148 24722 43204 24734
rect 43148 24670 43150 24722
rect 43202 24670 43204 24722
rect 43148 24164 43204 24670
rect 43148 24070 43204 24108
rect 43484 24724 43540 24734
rect 43484 24162 43540 24668
rect 43484 24110 43486 24162
rect 43538 24110 43540 24162
rect 43484 24098 43540 24110
rect 43372 23716 43428 23726
rect 43596 23716 43652 25230
rect 44716 24724 44772 24734
rect 44716 24630 44772 24668
rect 44380 24612 44436 24622
rect 44380 24518 44436 24556
rect 45164 23938 45220 25452
rect 45164 23886 45166 23938
rect 45218 23886 45220 23938
rect 45164 23874 45220 23886
rect 44828 23826 44884 23838
rect 44828 23774 44830 23826
rect 44882 23774 44884 23826
rect 43372 23714 43652 23716
rect 43372 23662 43374 23714
rect 43426 23662 43652 23714
rect 43372 23660 43652 23662
rect 44268 23714 44324 23726
rect 44268 23662 44270 23714
rect 44322 23662 44324 23714
rect 43148 23268 43204 23278
rect 43148 23042 43204 23212
rect 43148 22990 43150 23042
rect 43202 22990 43204 23042
rect 43036 22146 43092 22158
rect 43036 22094 43038 22146
rect 43090 22094 43092 22146
rect 43036 21924 43092 22094
rect 43036 21858 43092 21868
rect 42924 19292 43092 19348
rect 42588 18562 42644 18574
rect 42588 18510 42590 18562
rect 42642 18510 42644 18562
rect 42588 18452 42644 18510
rect 42588 18386 42644 18396
rect 42924 18450 42980 18462
rect 42924 18398 42926 18450
rect 42978 18398 42980 18450
rect 42924 18340 42980 18398
rect 42588 18228 42644 18238
rect 42588 17554 42644 18172
rect 42812 17892 42868 17902
rect 42812 17798 42868 17836
rect 42588 17502 42590 17554
rect 42642 17502 42644 17554
rect 42588 17490 42644 17502
rect 42700 17556 42756 17566
rect 42700 17462 42756 17500
rect 42812 17220 42868 17230
rect 42924 17220 42980 18284
rect 42476 17164 42644 17220
rect 42364 16716 42532 16772
rect 42364 16548 42420 16558
rect 42364 16322 42420 16492
rect 42364 16270 42366 16322
rect 42418 16270 42420 16322
rect 42364 16258 42420 16270
rect 42476 16212 42532 16716
rect 42476 16146 42532 16156
rect 42140 15932 42308 15988
rect 41916 14478 41918 14530
rect 41970 14478 41972 14530
rect 41916 14466 41972 14478
rect 42028 15428 42084 15438
rect 42028 15092 42084 15372
rect 42028 14308 42084 15036
rect 41804 13806 41806 13858
rect 41858 13806 41860 13858
rect 41804 13794 41860 13806
rect 41916 14252 42084 14308
rect 41692 13636 41748 13646
rect 41916 13636 41972 14252
rect 41692 13634 41972 13636
rect 41692 13582 41694 13634
rect 41746 13582 41972 13634
rect 41692 13580 41972 13582
rect 41692 13570 41748 13580
rect 42028 13524 42084 13534
rect 41916 13468 42028 13524
rect 41580 13074 41636 13086
rect 41580 13022 41582 13074
rect 41634 13022 41636 13074
rect 41468 12852 41524 12862
rect 41468 12758 41524 12796
rect 41244 10612 41300 10622
rect 41356 10612 41412 10780
rect 41244 10610 41412 10612
rect 41244 10558 41246 10610
rect 41298 10558 41412 10610
rect 41244 10556 41412 10558
rect 41468 10612 41524 10622
rect 41244 10546 41300 10556
rect 40908 10388 40964 10398
rect 40908 10386 41076 10388
rect 40908 10334 40910 10386
rect 40962 10334 41076 10386
rect 40908 10332 41076 10334
rect 40908 10322 40964 10332
rect 41020 10052 41076 10332
rect 41020 9714 41076 9996
rect 41020 9662 41022 9714
rect 41074 9662 41076 9714
rect 41020 9650 41076 9662
rect 41244 10386 41300 10398
rect 41244 10334 41246 10386
rect 41298 10334 41300 10386
rect 40684 9090 40740 9100
rect 41244 9042 41300 10334
rect 41468 9938 41524 10556
rect 41468 9886 41470 9938
rect 41522 9886 41524 9938
rect 41468 9874 41524 9886
rect 41244 8990 41246 9042
rect 41298 8990 41300 9042
rect 41244 8978 41300 8990
rect 41132 8932 41188 8942
rect 40572 8930 41188 8932
rect 40572 8878 41134 8930
rect 41186 8878 41188 8930
rect 40572 8876 41188 8878
rect 41132 8866 41188 8876
rect 41244 8820 41300 8830
rect 41244 8370 41300 8764
rect 41244 8318 41246 8370
rect 41298 8318 41300 8370
rect 41244 8306 41300 8318
rect 40572 8260 40628 8270
rect 40572 8166 40628 8204
rect 41132 7476 41188 7486
rect 41020 7474 41188 7476
rect 41020 7422 41134 7474
rect 41186 7422 41188 7474
rect 41020 7420 41188 7422
rect 40796 6804 40852 6814
rect 40460 6802 40852 6804
rect 40460 6750 40798 6802
rect 40850 6750 40852 6802
rect 40460 6748 40852 6750
rect 40796 6738 40852 6748
rect 40908 6692 40964 6702
rect 41020 6692 41076 7420
rect 41132 7410 41188 7420
rect 41580 7362 41636 13022
rect 41916 12850 41972 13468
rect 42028 13458 42084 13468
rect 41916 12798 41918 12850
rect 41970 12798 41972 12850
rect 41916 12786 41972 12798
rect 41692 12740 41748 12750
rect 41692 12646 41748 12684
rect 42028 12404 42084 12414
rect 42140 12404 42196 15932
rect 42476 15428 42532 15438
rect 42476 15314 42532 15372
rect 42476 15262 42478 15314
rect 42530 15262 42532 15314
rect 42476 15250 42532 15262
rect 42364 13076 42420 13086
rect 42364 12982 42420 13020
rect 42028 12402 42196 12404
rect 42028 12350 42030 12402
rect 42082 12350 42196 12402
rect 42028 12348 42196 12350
rect 42476 12516 42532 12526
rect 42028 12338 42084 12348
rect 42364 12068 42420 12078
rect 42252 11956 42308 11966
rect 42028 11900 42252 11956
rect 42028 11620 42084 11900
rect 42252 11890 42308 11900
rect 41916 11564 42084 11620
rect 41916 11170 41972 11564
rect 41916 11118 41918 11170
rect 41970 11118 41972 11170
rect 41916 11106 41972 11118
rect 42028 11394 42084 11406
rect 42028 11342 42030 11394
rect 42082 11342 42084 11394
rect 41692 10836 41748 10846
rect 41692 10742 41748 10780
rect 42028 10612 42084 11342
rect 42252 11396 42308 11406
rect 42364 11396 42420 12012
rect 42252 11394 42420 11396
rect 42252 11342 42254 11394
rect 42306 11342 42420 11394
rect 42252 11340 42420 11342
rect 42252 11330 42308 11340
rect 42028 10546 42084 10556
rect 42252 10500 42308 10510
rect 41804 10052 41860 10062
rect 41804 9826 41860 9996
rect 41804 9774 41806 9826
rect 41858 9774 41860 9826
rect 41804 9762 41860 9774
rect 42252 9826 42308 10444
rect 42364 10388 42420 11340
rect 42476 11284 42532 12460
rect 42588 11620 42644 17164
rect 42868 17164 42980 17220
rect 42812 17154 42868 17164
rect 43036 16100 43092 19292
rect 43036 16034 43092 16044
rect 42700 15876 42756 15886
rect 42700 15782 42756 15820
rect 42924 15316 42980 15326
rect 42924 15202 42980 15260
rect 42924 15150 42926 15202
rect 42978 15150 42980 15202
rect 42812 14308 42868 14318
rect 42812 13524 42868 14252
rect 42924 13636 42980 15150
rect 43148 15148 43204 22990
rect 43372 22148 43428 23660
rect 44268 23492 44324 23662
rect 44268 23426 44324 23436
rect 44380 23380 44436 23390
rect 44380 23378 44772 23380
rect 44380 23326 44382 23378
rect 44434 23326 44772 23378
rect 44380 23324 44772 23326
rect 44380 23314 44436 23324
rect 43372 22054 43428 22092
rect 43596 23156 43652 23166
rect 43596 21924 43652 23100
rect 44044 23154 44100 23166
rect 44044 23102 44046 23154
rect 44098 23102 44100 23154
rect 43596 21858 43652 21868
rect 43708 22484 43764 22494
rect 44044 22484 44100 23102
rect 44156 23156 44212 23166
rect 44156 23062 44212 23100
rect 44492 23154 44548 23166
rect 44492 23102 44494 23154
rect 44546 23102 44548 23154
rect 44492 22596 44548 23102
rect 44492 22530 44548 22540
rect 44044 22428 44324 22484
rect 43708 22370 43764 22428
rect 43708 22318 43710 22370
rect 43762 22318 43764 22370
rect 43484 21588 43540 21598
rect 43484 21494 43540 21532
rect 43708 21586 43764 22318
rect 43820 22372 43876 22382
rect 43820 22278 43876 22316
rect 43932 22148 43988 22158
rect 44156 22148 44212 22158
rect 43932 22054 43988 22092
rect 44044 22146 44212 22148
rect 44044 22094 44158 22146
rect 44210 22094 44212 22146
rect 44044 22092 44212 22094
rect 44044 21810 44100 22092
rect 44156 22082 44212 22092
rect 44044 21758 44046 21810
rect 44098 21758 44100 21810
rect 44044 21746 44100 21758
rect 44156 21924 44212 21934
rect 44156 21698 44212 21868
rect 44156 21646 44158 21698
rect 44210 21646 44212 21698
rect 44156 21634 44212 21646
rect 43708 21534 43710 21586
rect 43762 21534 43764 21586
rect 43708 21522 43764 21534
rect 44268 21588 44324 22428
rect 44716 22370 44772 23324
rect 44828 23266 44884 23774
rect 44828 23214 44830 23266
rect 44882 23214 44884 23266
rect 44828 23202 44884 23214
rect 44940 23716 44996 23726
rect 45276 23716 45332 27692
rect 45388 27682 45444 27692
rect 45612 27746 45892 27748
rect 45612 27694 45838 27746
rect 45890 27694 45892 27746
rect 45612 27692 45892 27694
rect 45612 27074 45668 27692
rect 45836 27682 45892 27692
rect 46396 27412 46452 27918
rect 54236 27970 54292 27982
rect 54236 27918 54238 27970
rect 54290 27918 54292 27970
rect 47292 27860 47348 27870
rect 46396 27346 46452 27356
rect 46732 27858 47348 27860
rect 46732 27806 47294 27858
rect 47346 27806 47348 27858
rect 46732 27804 47348 27806
rect 46732 27188 46788 27804
rect 47292 27794 47348 27804
rect 49644 27860 49700 27870
rect 47964 27748 48020 27758
rect 47964 27654 48020 27692
rect 49420 27746 49476 27758
rect 49420 27694 49422 27746
rect 49474 27694 49476 27746
rect 45612 27022 45614 27074
rect 45666 27022 45668 27074
rect 45612 26964 45668 27022
rect 46172 27132 46788 27188
rect 45612 26898 45668 26908
rect 45836 26964 45892 27002
rect 45836 26898 45892 26908
rect 46172 26850 46228 27132
rect 46508 26964 46564 26974
rect 46172 26798 46174 26850
rect 46226 26798 46228 26850
rect 46172 26740 46228 26798
rect 45724 26684 46228 26740
rect 46284 26850 46340 26862
rect 46284 26798 46286 26850
rect 46338 26798 46340 26850
rect 45724 26180 45780 26684
rect 46284 26628 46340 26798
rect 46396 26852 46452 26862
rect 46508 26852 46564 26908
rect 46396 26850 46564 26852
rect 46396 26798 46398 26850
rect 46450 26798 46564 26850
rect 46396 26796 46564 26798
rect 46396 26786 46452 26796
rect 45836 26572 46340 26628
rect 45836 26402 45892 26572
rect 46508 26514 46564 26796
rect 46508 26462 46510 26514
rect 46562 26462 46564 26514
rect 46508 26450 46564 26462
rect 45836 26350 45838 26402
rect 45890 26350 45892 26402
rect 45836 26338 45892 26350
rect 45948 26404 46004 26414
rect 46284 26404 46340 26414
rect 45948 26402 46340 26404
rect 45948 26350 45950 26402
rect 46002 26350 46286 26402
rect 46338 26350 46340 26402
rect 45948 26348 46340 26350
rect 45948 26338 46004 26348
rect 46284 26338 46340 26348
rect 46620 26404 46676 26414
rect 46732 26404 46788 27132
rect 46844 27412 46900 27422
rect 46844 27188 46900 27356
rect 47404 27412 47460 27422
rect 47404 27298 47460 27356
rect 49420 27412 49476 27694
rect 49420 27346 49476 27356
rect 49532 27748 49588 27758
rect 47404 27246 47406 27298
rect 47458 27246 47460 27298
rect 47404 27234 47460 27246
rect 49084 27300 49140 27338
rect 49084 27234 49140 27244
rect 46844 27132 47348 27188
rect 46844 27074 46900 27132
rect 46844 27022 46846 27074
rect 46898 27022 46900 27074
rect 46844 27010 46900 27022
rect 47068 26962 47124 26974
rect 47068 26910 47070 26962
rect 47122 26910 47124 26962
rect 47068 26908 47124 26910
rect 47292 26962 47348 27132
rect 49084 27074 49140 27086
rect 49084 27022 49086 27074
rect 49138 27022 49140 27074
rect 47292 26910 47294 26962
rect 47346 26910 47348 26962
rect 47292 26908 47348 26910
rect 46620 26402 46788 26404
rect 46620 26350 46622 26402
rect 46674 26350 46788 26402
rect 46620 26348 46788 26350
rect 46844 26852 47124 26908
rect 47180 26852 47348 26908
rect 48748 26964 48804 27002
rect 48748 26852 48916 26908
rect 46620 26338 46676 26348
rect 46508 26180 46564 26190
rect 45724 26124 45892 26180
rect 44940 23714 45332 23716
rect 44940 23662 44942 23714
rect 44994 23662 45332 23714
rect 44940 23660 45332 23662
rect 45612 24050 45668 24062
rect 45612 23998 45614 24050
rect 45666 23998 45668 24050
rect 44940 23492 44996 23660
rect 44716 22318 44718 22370
rect 44770 22318 44772 22370
rect 44716 22306 44772 22318
rect 44940 21924 44996 23436
rect 45388 23380 45444 23390
rect 45388 23154 45444 23324
rect 45388 23102 45390 23154
rect 45442 23102 45444 23154
rect 45388 23090 45444 23102
rect 45612 23042 45668 23998
rect 45612 22990 45614 23042
rect 45666 22990 45668 23042
rect 45388 22596 45444 22606
rect 45388 22482 45444 22540
rect 45388 22430 45390 22482
rect 45442 22430 45444 22482
rect 45388 22418 45444 22430
rect 45500 22370 45556 22382
rect 45500 22318 45502 22370
rect 45554 22318 45556 22370
rect 45500 22148 45556 22318
rect 45500 22082 45556 22092
rect 44940 21858 44996 21868
rect 44828 21812 44884 21822
rect 44828 21698 44884 21756
rect 44828 21646 44830 21698
rect 44882 21646 44884 21698
rect 44828 21634 44884 21646
rect 44380 21588 44436 21598
rect 44268 21586 44436 21588
rect 44268 21534 44382 21586
rect 44434 21534 44436 21586
rect 44268 21532 44436 21534
rect 44380 21364 44436 21532
rect 44716 21364 44772 21374
rect 44380 21362 44772 21364
rect 44380 21310 44718 21362
rect 44770 21310 44772 21362
rect 44380 21308 44772 21310
rect 44716 20580 44772 21308
rect 45388 20690 45444 20702
rect 45388 20638 45390 20690
rect 45442 20638 45444 20690
rect 44828 20580 44884 20590
rect 44716 20578 44884 20580
rect 44716 20526 44830 20578
rect 44882 20526 44884 20578
rect 44716 20524 44884 20526
rect 43932 19348 43988 19358
rect 43596 18676 43652 18686
rect 43372 18562 43428 18574
rect 43372 18510 43374 18562
rect 43426 18510 43428 18562
rect 43260 18450 43316 18462
rect 43260 18398 43262 18450
rect 43314 18398 43316 18450
rect 43260 17892 43316 18398
rect 43372 18452 43428 18510
rect 43372 18386 43428 18396
rect 43596 18450 43652 18620
rect 43596 18398 43598 18450
rect 43650 18398 43652 18450
rect 43596 18386 43652 18398
rect 43932 18450 43988 19292
rect 43932 18398 43934 18450
rect 43986 18398 43988 18450
rect 43932 18386 43988 18398
rect 44156 18450 44212 18462
rect 44156 18398 44158 18450
rect 44210 18398 44212 18450
rect 44156 18340 44212 18398
rect 44156 18274 44212 18284
rect 44604 18340 44660 18350
rect 43260 17826 43316 17836
rect 44604 16882 44660 18284
rect 44604 16830 44606 16882
rect 44658 16830 44660 16882
rect 44604 16818 44660 16830
rect 43596 16100 43652 16110
rect 43372 15988 43428 15998
rect 43372 15426 43428 15932
rect 43372 15374 43374 15426
rect 43426 15374 43428 15426
rect 43372 15362 43428 15374
rect 43148 15092 43316 15148
rect 43148 14420 43204 14430
rect 43148 14326 43204 14364
rect 43036 13746 43092 13758
rect 43036 13694 43038 13746
rect 43090 13694 43092 13746
rect 43036 13636 43092 13694
rect 42980 13580 43092 13636
rect 42924 13570 42980 13580
rect 42812 13458 42868 13468
rect 43148 12962 43204 12974
rect 43148 12910 43150 12962
rect 43202 12910 43204 12962
rect 42924 12178 42980 12190
rect 42924 12126 42926 12178
rect 42978 12126 42980 12178
rect 42812 12068 42868 12078
rect 42924 12068 42980 12126
rect 42868 12012 42980 12068
rect 42812 12002 42868 12012
rect 43148 11956 43204 12910
rect 43148 11890 43204 11900
rect 42812 11620 42868 11630
rect 42588 11618 42868 11620
rect 42588 11566 42814 11618
rect 42866 11566 42868 11618
rect 42588 11564 42868 11566
rect 42588 11284 42644 11294
rect 42476 11282 42756 11284
rect 42476 11230 42590 11282
rect 42642 11230 42756 11282
rect 42476 11228 42756 11230
rect 42588 11218 42644 11228
rect 42700 10836 42756 11228
rect 42812 11060 42868 11564
rect 43260 11508 43316 15092
rect 43596 14642 43652 16044
rect 43932 16100 43988 16110
rect 43932 16006 43988 16044
rect 44156 16100 44212 16110
rect 44156 15986 44212 16044
rect 44156 15934 44158 15986
rect 44210 15934 44212 15986
rect 44156 15922 44212 15934
rect 44716 15148 44772 20524
rect 44828 20514 44884 20524
rect 45388 20580 45444 20638
rect 45276 20020 45332 20030
rect 44828 18564 44884 18574
rect 44828 18450 44884 18508
rect 44828 18398 44830 18450
rect 44882 18398 44884 18450
rect 44828 18386 44884 18398
rect 45164 17556 45220 17566
rect 45164 17462 45220 17500
rect 45052 16994 45108 17006
rect 45052 16942 45054 16994
rect 45106 16942 45108 16994
rect 45052 16772 45108 16942
rect 45052 16100 45108 16716
rect 45276 16770 45332 19964
rect 45388 17444 45444 20524
rect 45500 20020 45556 20030
rect 45612 20020 45668 22990
rect 45556 19964 45668 20020
rect 45500 19954 45556 19964
rect 45724 18676 45780 18686
rect 45724 18562 45780 18620
rect 45724 18510 45726 18562
rect 45778 18510 45780 18562
rect 45724 18498 45780 18510
rect 45612 18452 45668 18462
rect 45500 18450 45668 18452
rect 45500 18398 45614 18450
rect 45666 18398 45668 18450
rect 45500 18396 45668 18398
rect 45500 17890 45556 18396
rect 45612 18386 45668 18396
rect 45836 18338 45892 26124
rect 45948 26066 46004 26078
rect 45948 26014 45950 26066
rect 46002 26014 46004 26066
rect 45948 24948 46004 26014
rect 46284 25508 46340 25518
rect 46284 25414 46340 25452
rect 46508 25506 46564 26124
rect 46508 25454 46510 25506
rect 46562 25454 46564 25506
rect 46508 25284 46564 25454
rect 46844 25508 46900 26852
rect 47068 26516 47124 26526
rect 47180 26516 47236 26852
rect 47068 26514 47236 26516
rect 47068 26462 47070 26514
rect 47122 26462 47236 26514
rect 47068 26460 47236 26462
rect 47068 26450 47124 26460
rect 48860 26290 48916 26852
rect 48860 26238 48862 26290
rect 48914 26238 48916 26290
rect 48860 26226 48916 26238
rect 49084 26290 49140 27022
rect 49532 27074 49588 27692
rect 49644 27300 49700 27804
rect 50428 27858 50484 27870
rect 50428 27806 50430 27858
rect 50482 27806 50484 27858
rect 49868 27748 49924 27758
rect 49868 27654 49924 27692
rect 50428 27748 50484 27806
rect 50428 27682 50484 27692
rect 50876 27858 50932 27870
rect 50876 27806 50878 27858
rect 50930 27806 50932 27858
rect 50316 27636 50372 27646
rect 50316 27542 50372 27580
rect 49980 27412 50036 27422
rect 49756 27300 49812 27310
rect 49700 27298 49812 27300
rect 49700 27246 49758 27298
rect 49810 27246 49812 27298
rect 49700 27244 49812 27246
rect 49644 27206 49700 27244
rect 49756 27234 49812 27244
rect 49980 27298 50036 27356
rect 50876 27412 50932 27806
rect 51100 27860 51156 27870
rect 51100 27766 51156 27804
rect 51996 27860 52052 27870
rect 50988 27746 51044 27758
rect 50988 27694 50990 27746
rect 51042 27694 51044 27746
rect 50988 27636 51044 27694
rect 51436 27746 51492 27758
rect 51436 27694 51438 27746
rect 51490 27694 51492 27746
rect 51436 27636 51492 27694
rect 50988 27580 51492 27636
rect 51436 27412 51492 27580
rect 51660 27636 51716 27646
rect 51660 27542 51716 27580
rect 51436 27356 51940 27412
rect 50876 27346 50932 27356
rect 49980 27246 49982 27298
rect 50034 27246 50036 27298
rect 49980 27234 50036 27246
rect 49532 27022 49534 27074
rect 49586 27022 49588 27074
rect 49532 27010 49588 27022
rect 51772 27076 51828 27086
rect 51772 26982 51828 27020
rect 50092 26962 50148 26974
rect 50092 26910 50094 26962
rect 50146 26910 50148 26962
rect 49756 26404 49812 26414
rect 49756 26310 49812 26348
rect 49084 26238 49086 26290
rect 49138 26238 49140 26290
rect 46956 26180 47012 26190
rect 46956 26086 47012 26124
rect 47180 25620 47236 25630
rect 47180 25526 47236 25564
rect 49084 25620 49140 26238
rect 50092 26292 50148 26910
rect 50876 26964 50932 26974
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50316 26404 50372 26414
rect 50372 26348 50484 26404
rect 50316 26310 50372 26348
rect 50092 26226 50148 26236
rect 50204 26290 50260 26302
rect 50204 26238 50206 26290
rect 50258 26238 50260 26290
rect 49084 25554 49140 25564
rect 46844 25442 46900 25452
rect 48860 25508 48916 25518
rect 46508 25218 46564 25228
rect 46956 25284 47012 25294
rect 45948 24892 46788 24948
rect 46284 24724 46340 24734
rect 46060 23938 46116 23950
rect 46060 23886 46062 23938
rect 46114 23886 46116 23938
rect 46060 22036 46116 23886
rect 46060 21970 46116 21980
rect 46172 22258 46228 22270
rect 46172 22206 46174 22258
rect 46226 22206 46228 22258
rect 45836 18286 45838 18338
rect 45890 18286 45892 18338
rect 45836 18274 45892 18286
rect 45948 21924 46004 21934
rect 45500 17838 45502 17890
rect 45554 17838 45556 17890
rect 45500 17826 45556 17838
rect 45500 17668 45556 17678
rect 45500 17574 45556 17612
rect 45388 17388 45668 17444
rect 45276 16718 45278 16770
rect 45330 16718 45332 16770
rect 45276 16706 45332 16718
rect 45500 16882 45556 16894
rect 45500 16830 45502 16882
rect 45554 16830 45556 16882
rect 45500 16772 45556 16830
rect 45164 16324 45220 16334
rect 45500 16324 45556 16716
rect 45164 16322 45556 16324
rect 45164 16270 45166 16322
rect 45218 16270 45556 16322
rect 45164 16268 45556 16270
rect 45164 16258 45220 16268
rect 45164 16100 45220 16110
rect 45052 16098 45220 16100
rect 45052 16046 45166 16098
rect 45218 16046 45220 16098
rect 45052 16044 45220 16046
rect 44828 15988 44884 15998
rect 44828 15894 44884 15932
rect 45164 15764 45220 16044
rect 45164 15698 45220 15708
rect 43596 14590 43598 14642
rect 43650 14590 43652 14642
rect 43596 14578 43652 14590
rect 44156 15092 44772 15148
rect 45612 15148 45668 17388
rect 45948 15202 46004 21868
rect 46172 21364 46228 22206
rect 46172 21298 46228 21308
rect 46172 20580 46228 20590
rect 46284 20580 46340 24668
rect 46732 23938 46788 24892
rect 46844 24164 46900 24174
rect 46844 24070 46900 24108
rect 46956 24050 47012 25228
rect 48860 24946 48916 25452
rect 50204 25508 50260 26238
rect 50428 25956 50484 26348
rect 50540 26292 50596 26302
rect 50764 26292 50820 26302
rect 50876 26292 50932 26908
rect 51436 26962 51492 26974
rect 51436 26910 51438 26962
rect 51490 26910 51492 26962
rect 50540 26290 50932 26292
rect 50540 26238 50542 26290
rect 50594 26238 50766 26290
rect 50818 26238 50932 26290
rect 50540 26236 50932 26238
rect 50988 26292 51044 26302
rect 50540 26226 50596 26236
rect 50764 26226 50820 26236
rect 50988 26198 51044 26236
rect 51436 26292 51492 26910
rect 51436 26226 51492 26236
rect 51660 26962 51716 26974
rect 51660 26910 51662 26962
rect 51714 26910 51716 26962
rect 50764 26066 50820 26078
rect 50764 26014 50766 26066
rect 50818 26014 50820 26066
rect 50540 25956 50596 25966
rect 50428 25900 50540 25956
rect 50540 25890 50596 25900
rect 50204 25442 50260 25452
rect 50652 25508 50708 25518
rect 50652 25414 50708 25452
rect 50764 25284 50820 26014
rect 50876 25956 50932 25966
rect 50876 25506 50932 25900
rect 51548 25620 51604 25630
rect 51660 25620 51716 26910
rect 51884 26908 51940 27356
rect 51996 27076 52052 27804
rect 52892 27860 52948 27870
rect 52892 27766 52948 27804
rect 53564 27860 53620 27870
rect 53900 27860 53956 27870
rect 53564 27858 53956 27860
rect 53564 27806 53566 27858
rect 53618 27806 53902 27858
rect 53954 27806 53956 27858
rect 53564 27804 53956 27806
rect 53564 27794 53620 27804
rect 53900 27794 53956 27804
rect 53116 27746 53172 27758
rect 53116 27694 53118 27746
rect 53170 27694 53172 27746
rect 53116 27186 53172 27694
rect 53116 27134 53118 27186
rect 53170 27134 53172 27186
rect 53116 27122 53172 27134
rect 51996 27010 52052 27020
rect 52556 27074 52612 27086
rect 52556 27022 52558 27074
rect 52610 27022 52612 27074
rect 52556 26964 52612 27022
rect 54236 27076 54292 27918
rect 57932 27636 57988 27646
rect 57932 27298 57988 27580
rect 57932 27246 57934 27298
rect 57986 27246 57988 27298
rect 57932 27234 57988 27246
rect 54236 27010 54292 27020
rect 55580 27076 55636 27086
rect 55580 26982 55636 27020
rect 51884 26852 52052 26908
rect 52556 26898 52612 26908
rect 53004 26852 53060 26862
rect 51996 26290 52052 26852
rect 52892 26850 53060 26852
rect 52892 26798 53006 26850
rect 53058 26798 53060 26850
rect 52892 26796 53060 26798
rect 51996 26238 51998 26290
rect 52050 26238 52052 26290
rect 51996 26226 52052 26238
rect 52332 26292 52388 26302
rect 52332 26198 52388 26236
rect 52892 26292 52948 26796
rect 53004 26786 53060 26796
rect 53228 26850 53284 26862
rect 53228 26798 53230 26850
rect 53282 26798 53284 26850
rect 52780 25732 52836 25742
rect 52892 25732 52948 26236
rect 53004 26290 53060 26302
rect 53004 26238 53006 26290
rect 53058 26238 53060 26290
rect 53004 26180 53060 26238
rect 53228 26180 53284 26798
rect 55020 26402 55076 26414
rect 55020 26350 55022 26402
rect 55074 26350 55076 26402
rect 53676 26292 53732 26302
rect 53676 26198 53732 26236
rect 54348 26292 54404 26302
rect 54684 26292 54740 26302
rect 54348 26290 54740 26292
rect 54348 26238 54350 26290
rect 54402 26238 54686 26290
rect 54738 26238 54740 26290
rect 54348 26236 54740 26238
rect 54348 26226 54404 26236
rect 54684 26226 54740 26236
rect 53564 26180 53620 26190
rect 53004 26178 53620 26180
rect 53004 26126 53566 26178
rect 53618 26126 53620 26178
rect 53004 26124 53620 26126
rect 53564 26068 53620 26124
rect 53564 26012 53732 26068
rect 52780 25730 52948 25732
rect 52780 25678 52782 25730
rect 52834 25678 52948 25730
rect 52780 25676 52948 25678
rect 52780 25666 52836 25676
rect 51548 25618 51660 25620
rect 51548 25566 51550 25618
rect 51602 25566 51660 25618
rect 51548 25564 51660 25566
rect 51548 25554 51604 25564
rect 51660 25526 51716 25564
rect 52668 25620 52724 25630
rect 52668 25526 52724 25564
rect 50876 25454 50878 25506
rect 50930 25454 50932 25506
rect 50876 25442 50932 25454
rect 50764 25218 50820 25228
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 53004 24948 53060 24958
rect 48860 24894 48862 24946
rect 48914 24894 48916 24946
rect 48860 24882 48916 24894
rect 49084 24892 49588 24948
rect 47068 24724 47124 24734
rect 47068 24630 47124 24668
rect 47964 24724 48020 24734
rect 46956 23998 46958 24050
rect 47010 23998 47012 24050
rect 46956 23986 47012 23998
rect 46732 23886 46734 23938
rect 46786 23886 46788 23938
rect 46732 23874 46788 23886
rect 47180 23940 47236 23950
rect 46732 21700 46788 21710
rect 46620 21698 46788 21700
rect 46620 21646 46734 21698
rect 46786 21646 46788 21698
rect 46620 21644 46788 21646
rect 46228 20524 46340 20580
rect 46396 20802 46452 20814
rect 46396 20750 46398 20802
rect 46450 20750 46452 20802
rect 46396 20692 46452 20750
rect 46172 20514 46228 20524
rect 46172 19348 46228 19358
rect 46396 19348 46452 20636
rect 46620 20802 46676 21644
rect 46732 21634 46788 21644
rect 46844 21588 46900 21598
rect 47068 21588 47124 21598
rect 46844 21494 46900 21532
rect 46956 21586 47124 21588
rect 46956 21534 47070 21586
rect 47122 21534 47124 21586
rect 46956 21532 47124 21534
rect 46732 21364 46788 21374
rect 46956 21364 47012 21532
rect 47068 21522 47124 21532
rect 46732 21362 47012 21364
rect 46732 21310 46734 21362
rect 46786 21310 47012 21362
rect 46732 21308 47012 21310
rect 46732 21298 46788 21308
rect 46620 20750 46622 20802
rect 46674 20750 46676 20802
rect 46620 20244 46676 20750
rect 46620 20178 46676 20188
rect 46172 19346 46452 19348
rect 46172 19294 46174 19346
rect 46226 19294 46452 19346
rect 46172 19292 46452 19294
rect 46844 20132 46900 20142
rect 46172 19282 46228 19292
rect 46620 19236 46676 19246
rect 46620 19142 46676 19180
rect 46060 19012 46116 19022
rect 46060 18918 46116 18956
rect 46284 19012 46340 19022
rect 46284 18918 46340 18956
rect 46620 18450 46676 18462
rect 46620 18398 46622 18450
rect 46674 18398 46676 18450
rect 46396 17666 46452 17678
rect 46396 17614 46398 17666
rect 46450 17614 46452 17666
rect 46284 16996 46340 17006
rect 46172 16994 46340 16996
rect 46172 16942 46286 16994
rect 46338 16942 46340 16994
rect 46172 16940 46340 16942
rect 46060 16772 46116 16782
rect 46060 16678 46116 16716
rect 45948 15150 45950 15202
rect 46002 15150 46004 15202
rect 45612 15092 45780 15148
rect 43484 14308 43540 14318
rect 43484 14214 43540 14252
rect 43484 13970 43540 13982
rect 43484 13918 43486 13970
rect 43538 13918 43540 13970
rect 43372 13074 43428 13086
rect 43372 13022 43374 13074
rect 43426 13022 43428 13074
rect 43372 12964 43428 13022
rect 43372 12898 43428 12908
rect 43260 11442 43316 11452
rect 43372 11394 43428 11406
rect 43372 11342 43374 11394
rect 43426 11342 43428 11394
rect 43372 11172 43428 11342
rect 42812 10994 42868 11004
rect 42924 11116 43428 11172
rect 42812 10836 42868 10846
rect 42700 10834 42868 10836
rect 42700 10782 42814 10834
rect 42866 10782 42868 10834
rect 42700 10780 42868 10782
rect 42812 10770 42868 10780
rect 42812 10500 42868 10510
rect 42700 10444 42812 10500
rect 42588 10388 42644 10398
rect 42364 10386 42644 10388
rect 42364 10334 42590 10386
rect 42642 10334 42644 10386
rect 42364 10332 42644 10334
rect 42252 9774 42254 9826
rect 42306 9774 42308 9826
rect 42252 9762 42308 9774
rect 41580 7310 41582 7362
rect 41634 7310 41636 7362
rect 41580 7298 41636 7310
rect 41692 9714 41748 9726
rect 41692 9662 41694 9714
rect 41746 9662 41748 9714
rect 40964 6636 41076 6692
rect 41356 6692 41412 6702
rect 40908 6598 40964 6636
rect 41356 6598 41412 6636
rect 40348 6402 40404 6412
rect 41692 6356 41748 9662
rect 42588 9604 42644 10332
rect 42140 9548 42644 9604
rect 42028 9156 42084 9166
rect 42028 9062 42084 9100
rect 41916 7252 41972 7262
rect 41972 7196 42084 7252
rect 41916 7158 41972 7196
rect 41916 6580 41972 6590
rect 41916 6486 41972 6524
rect 40236 5966 40238 6018
rect 40290 5966 40292 6018
rect 40236 5954 40292 5966
rect 41244 6300 41748 6356
rect 39788 5908 39844 5918
rect 40124 5908 40180 5918
rect 39340 5906 40180 5908
rect 39340 5854 39790 5906
rect 39842 5854 40126 5906
rect 40178 5854 40180 5906
rect 39340 5852 40180 5854
rect 39340 5122 39396 5852
rect 39788 5842 39844 5852
rect 40124 5842 40180 5852
rect 39452 5684 39508 5694
rect 39452 5590 39508 5628
rect 39788 5684 39844 5694
rect 39788 5682 40068 5684
rect 39788 5630 39790 5682
rect 39842 5630 40068 5682
rect 39788 5628 40068 5630
rect 39788 5618 39844 5628
rect 39340 5070 39342 5122
rect 39394 5070 39396 5122
rect 39340 5058 39396 5070
rect 39788 5124 39844 5134
rect 40012 5124 40068 5628
rect 41132 5236 41188 5246
rect 41132 5142 41188 5180
rect 40124 5124 40180 5134
rect 40012 5122 40180 5124
rect 40012 5070 40126 5122
rect 40178 5070 40180 5122
rect 40012 5068 40180 5070
rect 39676 5012 39732 5022
rect 39676 4338 39732 4956
rect 39676 4286 39678 4338
rect 39730 4286 39732 4338
rect 39676 4274 39732 4286
rect 39788 4228 39844 5068
rect 40124 5058 40180 5068
rect 40684 5124 40740 5134
rect 40684 5030 40740 5068
rect 41244 5012 41300 6300
rect 42028 5906 42084 7196
rect 42140 6020 42196 9548
rect 42700 8932 42756 10444
rect 42812 10434 42868 10444
rect 42924 10498 42980 11116
rect 43372 10948 43428 10958
rect 43372 10834 43428 10892
rect 43372 10782 43374 10834
rect 43426 10782 43428 10834
rect 43372 10770 43428 10782
rect 43260 10612 43316 10622
rect 43260 10518 43316 10556
rect 42924 10446 42926 10498
rect 42978 10446 42980 10498
rect 42924 10434 42980 10446
rect 43484 10052 43540 13918
rect 43932 12964 43988 12974
rect 43820 12850 43876 12862
rect 43820 12798 43822 12850
rect 43874 12798 43876 12850
rect 43820 12180 43876 12798
rect 43932 12290 43988 12908
rect 43932 12238 43934 12290
rect 43986 12238 43988 12290
rect 43932 12226 43988 12238
rect 43820 12114 43876 12124
rect 43596 11506 43652 11518
rect 43596 11454 43598 11506
rect 43650 11454 43652 11506
rect 43596 10834 43652 11454
rect 43596 10782 43598 10834
rect 43650 10782 43652 10834
rect 43596 10770 43652 10782
rect 43484 9986 43540 9996
rect 42812 9714 42868 9726
rect 42812 9662 42814 9714
rect 42866 9662 42868 9714
rect 42812 9156 42868 9662
rect 42924 9604 42980 9614
rect 43148 9604 43204 9614
rect 42924 9510 42980 9548
rect 43036 9602 43204 9604
rect 43036 9550 43150 9602
rect 43202 9550 43204 9602
rect 43036 9548 43204 9550
rect 42812 9090 42868 9100
rect 42812 8932 42868 8942
rect 42700 8930 42868 8932
rect 42700 8878 42814 8930
rect 42866 8878 42868 8930
rect 42700 8876 42868 8878
rect 42812 8866 42868 8876
rect 43036 7364 43092 9548
rect 43148 9538 43204 9548
rect 43484 9604 43540 9614
rect 43484 9510 43540 9548
rect 44156 9266 44212 15092
rect 45500 14642 45556 14654
rect 45500 14590 45502 14642
rect 45554 14590 45556 14642
rect 45388 14530 45444 14542
rect 45388 14478 45390 14530
rect 45442 14478 45444 14530
rect 45388 13748 45444 14478
rect 45388 13654 45444 13692
rect 45500 14532 45556 14590
rect 45500 13636 45556 14476
rect 45612 13636 45668 13646
rect 45500 13634 45668 13636
rect 45500 13582 45614 13634
rect 45666 13582 45668 13634
rect 45500 13580 45668 13582
rect 45612 13570 45668 13580
rect 44268 12964 44324 12974
rect 44268 12870 44324 12908
rect 45052 12180 45108 12190
rect 44940 12178 45108 12180
rect 44940 12126 45054 12178
rect 45106 12126 45108 12178
rect 44940 12124 45108 12126
rect 44268 11284 44324 11294
rect 44268 11282 44884 11284
rect 44268 11230 44270 11282
rect 44322 11230 44884 11282
rect 44268 11228 44884 11230
rect 44268 11218 44324 11228
rect 44828 10610 44884 11228
rect 44828 10558 44830 10610
rect 44882 10558 44884 10610
rect 44828 10546 44884 10558
rect 44940 10612 44996 12124
rect 45052 12114 45108 12124
rect 45388 12180 45444 12190
rect 45388 12086 45444 12124
rect 45724 12178 45780 15092
rect 45948 14868 46004 15150
rect 46172 16100 46228 16940
rect 46284 16930 46340 16940
rect 46396 16770 46452 17614
rect 46396 16718 46398 16770
rect 46450 16718 46452 16770
rect 46396 16706 46452 16718
rect 46172 15148 46228 16044
rect 45948 14802 46004 14812
rect 46060 15092 46228 15148
rect 46508 15764 46564 15774
rect 46060 14644 46116 15092
rect 46508 14868 46564 15708
rect 46620 15148 46676 18398
rect 46844 17778 46900 20076
rect 46956 19908 47012 19918
rect 46956 19234 47012 19852
rect 47068 19348 47124 19358
rect 47180 19348 47236 23884
rect 47964 23938 48020 24668
rect 48748 24722 48804 24734
rect 48748 24670 48750 24722
rect 48802 24670 48804 24722
rect 47964 23886 47966 23938
rect 48018 23886 48020 23938
rect 47964 23604 48020 23886
rect 48188 24050 48244 24062
rect 48188 23998 48190 24050
rect 48242 23998 48244 24050
rect 48188 23940 48244 23998
rect 48188 23874 48244 23884
rect 48748 23940 48804 24670
rect 48972 24724 49028 24734
rect 48972 24630 49028 24668
rect 49084 24276 49140 24892
rect 49532 24836 49588 24892
rect 52780 24946 53060 24948
rect 52780 24894 53006 24946
rect 53058 24894 53060 24946
rect 52780 24892 53060 24894
rect 49644 24836 49700 24846
rect 49532 24834 49700 24836
rect 49532 24782 49646 24834
rect 49698 24782 49700 24834
rect 49532 24780 49700 24782
rect 49644 24770 49700 24780
rect 49420 24722 49476 24734
rect 49420 24670 49422 24722
rect 49474 24670 49476 24722
rect 48748 23874 48804 23884
rect 48860 24220 49140 24276
rect 49308 24612 49364 24622
rect 48860 23938 48916 24220
rect 49308 24052 49364 24556
rect 48860 23886 48862 23938
rect 48914 23886 48916 23938
rect 48860 23874 48916 23886
rect 49196 24050 49364 24052
rect 49196 23998 49310 24050
rect 49362 23998 49364 24050
rect 49196 23996 49364 23998
rect 47964 23538 48020 23548
rect 47628 23268 47684 23278
rect 47292 23044 47348 23054
rect 47292 22484 47348 22988
rect 47292 22390 47348 22428
rect 47404 23042 47460 23054
rect 47404 22990 47406 23042
rect 47458 22990 47460 23042
rect 47404 22036 47460 22990
rect 47404 21970 47460 21980
rect 47516 22370 47572 22382
rect 47516 22318 47518 22370
rect 47570 22318 47572 22370
rect 47516 21812 47572 22318
rect 47292 21810 47572 21812
rect 47292 21758 47518 21810
rect 47570 21758 47572 21810
rect 47292 21756 47572 21758
rect 47292 20914 47348 21756
rect 47516 21746 47572 21756
rect 47628 21810 47684 23212
rect 49196 23266 49252 23996
rect 49308 23986 49364 23996
rect 49420 23380 49476 24670
rect 49756 24498 49812 24510
rect 49756 24446 49758 24498
rect 49810 24446 49812 24498
rect 49756 23938 49812 24446
rect 49756 23886 49758 23938
rect 49810 23886 49812 23938
rect 49532 23380 49588 23390
rect 49420 23378 49588 23380
rect 49420 23326 49534 23378
rect 49586 23326 49588 23378
rect 49420 23324 49588 23326
rect 49532 23314 49588 23324
rect 49196 23214 49198 23266
rect 49250 23214 49252 23266
rect 49196 23202 49252 23214
rect 49308 23266 49364 23278
rect 49308 23214 49310 23266
rect 49362 23214 49364 23266
rect 49308 23156 49364 23214
rect 49756 23156 49812 23886
rect 50204 23826 50260 23838
rect 50204 23774 50206 23826
rect 50258 23774 50260 23826
rect 50204 23380 50260 23774
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 51436 23492 51492 23502
rect 50204 23314 50260 23324
rect 51100 23380 51156 23390
rect 51100 23266 51156 23324
rect 51436 23378 51492 23436
rect 52780 23492 52836 24892
rect 53004 24882 53060 24892
rect 51436 23326 51438 23378
rect 51490 23326 51492 23378
rect 51436 23314 51492 23326
rect 51884 23380 51940 23390
rect 51100 23214 51102 23266
rect 51154 23214 51156 23266
rect 51100 23202 51156 23214
rect 51212 23268 51268 23278
rect 51212 23174 51268 23212
rect 51660 23268 51716 23278
rect 51660 23174 51716 23212
rect 49308 23100 49812 23156
rect 51884 23154 51940 23324
rect 52220 23380 52276 23390
rect 52220 23286 52276 23324
rect 52668 23380 52724 23390
rect 52780 23380 52836 23436
rect 52668 23378 52836 23380
rect 52668 23326 52670 23378
rect 52722 23326 52836 23378
rect 52668 23324 52836 23326
rect 52892 24722 52948 24734
rect 52892 24670 52894 24722
rect 52946 24670 52948 24722
rect 52892 23938 52948 24670
rect 53228 24722 53284 24734
rect 53228 24670 53230 24722
rect 53282 24670 53284 24722
rect 53228 24276 53284 24670
rect 53228 24220 53620 24276
rect 53340 24052 53396 24062
rect 52892 23886 52894 23938
rect 52946 23886 52948 23938
rect 52892 23380 52948 23886
rect 52668 23314 52724 23324
rect 52892 23314 52948 23324
rect 53004 24050 53396 24052
rect 53004 23998 53342 24050
rect 53394 23998 53396 24050
rect 53004 23996 53396 23998
rect 53004 23378 53060 23996
rect 53340 23986 53396 23996
rect 53004 23326 53006 23378
rect 53058 23326 53060 23378
rect 53004 23314 53060 23326
rect 53452 23938 53508 23950
rect 53452 23886 53454 23938
rect 53506 23886 53508 23938
rect 51884 23102 51886 23154
rect 51938 23102 51940 23154
rect 51884 23090 51940 23102
rect 52892 23154 52948 23166
rect 52892 23102 52894 23154
rect 52946 23102 52948 23154
rect 52892 22708 52948 23102
rect 53116 23156 53172 23166
rect 53116 23154 53284 23156
rect 53116 23102 53118 23154
rect 53170 23102 53284 23154
rect 53116 23100 53284 23102
rect 53116 23090 53172 23100
rect 50764 22652 51044 22708
rect 47964 22596 48020 22606
rect 47964 22502 48020 22540
rect 50764 22594 50820 22652
rect 50764 22542 50766 22594
rect 50818 22542 50820 22594
rect 50764 22530 50820 22542
rect 47628 21758 47630 21810
rect 47682 21758 47684 21810
rect 47628 21746 47684 21758
rect 47740 22484 47796 22494
rect 47740 21810 47796 22428
rect 50876 22484 50932 22494
rect 50204 22372 50260 22382
rect 50204 22278 50260 22316
rect 50428 22370 50484 22382
rect 50428 22318 50430 22370
rect 50482 22318 50484 22370
rect 50428 21924 50484 22318
rect 50652 22370 50708 22382
rect 50652 22318 50654 22370
rect 50706 22318 50708 22370
rect 50652 22148 50708 22318
rect 50652 22082 50708 22092
rect 47740 21758 47742 21810
rect 47794 21758 47796 21810
rect 47740 21746 47796 21758
rect 49980 21868 50484 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 49420 21700 49476 21710
rect 47404 21588 47460 21598
rect 47460 21532 47572 21588
rect 47404 21522 47460 21532
rect 47516 21028 47572 21532
rect 49196 21140 49252 21150
rect 47628 21028 47684 21038
rect 47516 21026 47684 21028
rect 47516 20974 47630 21026
rect 47682 20974 47684 21026
rect 47516 20972 47684 20974
rect 47628 20962 47684 20972
rect 47292 20862 47294 20914
rect 47346 20862 47348 20914
rect 47292 20850 47348 20862
rect 47740 20692 47796 20702
rect 47740 20598 47796 20636
rect 47068 19346 47236 19348
rect 47068 19294 47070 19346
rect 47122 19294 47236 19346
rect 47068 19292 47236 19294
rect 47068 19282 47124 19292
rect 46956 19182 46958 19234
rect 47010 19182 47012 19234
rect 46956 19170 47012 19182
rect 47628 19236 47684 19246
rect 46956 19012 47012 19022
rect 47180 19012 47236 19022
rect 47012 19010 47236 19012
rect 47012 18958 47182 19010
rect 47234 18958 47236 19010
rect 47012 18956 47236 18958
rect 46956 18340 47012 18956
rect 47180 18946 47236 18956
rect 47068 18564 47124 18574
rect 47068 18470 47124 18508
rect 47180 18452 47236 18462
rect 47180 18358 47236 18396
rect 47292 18452 47348 18462
rect 47628 18452 47684 19180
rect 47740 18452 47796 18462
rect 47292 18450 47460 18452
rect 47292 18398 47294 18450
rect 47346 18398 47460 18450
rect 47292 18396 47460 18398
rect 47628 18450 47796 18452
rect 47628 18398 47742 18450
rect 47794 18398 47796 18450
rect 47628 18396 47796 18398
rect 47292 18386 47348 18396
rect 46956 18284 47124 18340
rect 46844 17726 46846 17778
rect 46898 17726 46900 17778
rect 46844 17714 46900 17726
rect 47068 17668 47124 18284
rect 46732 17442 46788 17454
rect 46732 17390 46734 17442
rect 46786 17390 46788 17442
rect 46732 17108 46788 17390
rect 46956 17444 47012 17454
rect 47068 17444 47124 17612
rect 47292 17444 47348 17454
rect 47068 17442 47348 17444
rect 47068 17390 47294 17442
rect 47346 17390 47348 17442
rect 47068 17388 47348 17390
rect 47404 17444 47460 18396
rect 47628 17444 47684 17454
rect 47404 17388 47628 17444
rect 46956 17350 47012 17388
rect 47292 17332 47348 17388
rect 47628 17350 47684 17388
rect 47292 17276 47460 17332
rect 47068 17108 47124 17118
rect 46732 17052 47068 17108
rect 47068 17014 47124 17052
rect 46732 16882 46788 16894
rect 46732 16830 46734 16882
rect 46786 16830 46788 16882
rect 46732 15876 46788 16830
rect 47180 16210 47236 16222
rect 47180 16158 47182 16210
rect 47234 16158 47236 16210
rect 46732 15810 46788 15820
rect 46956 16098 47012 16110
rect 46956 16046 46958 16098
rect 47010 16046 47012 16098
rect 46956 15148 47012 16046
rect 47180 16100 47236 16158
rect 47180 16034 47236 16044
rect 47068 15986 47124 15998
rect 47068 15934 47070 15986
rect 47122 15934 47124 15986
rect 47068 15876 47124 15934
rect 47068 15810 47124 15820
rect 46620 15092 46900 15148
rect 46956 15092 47236 15148
rect 46508 14802 46564 14812
rect 45724 12126 45726 12178
rect 45778 12126 45780 12178
rect 44940 10546 44996 10556
rect 45164 11508 45220 11518
rect 45164 10610 45220 11452
rect 45164 10558 45166 10610
rect 45218 10558 45220 10610
rect 45164 10500 45220 10558
rect 45164 10434 45220 10444
rect 45724 11508 45780 12126
rect 45052 10388 45108 10398
rect 44156 9214 44158 9266
rect 44210 9214 44212 9266
rect 44156 9202 44212 9214
rect 44604 10052 44660 10062
rect 44604 9154 44660 9996
rect 44604 9102 44606 9154
rect 44658 9102 44660 9154
rect 44604 8932 44660 9102
rect 44828 9156 44884 9166
rect 45052 9156 45108 10332
rect 45500 10386 45556 10398
rect 45500 10334 45502 10386
rect 45554 10334 45556 10386
rect 44828 9154 45108 9156
rect 44828 9102 44830 9154
rect 44882 9102 45108 9154
rect 44828 9100 45108 9102
rect 45276 9268 45332 9278
rect 44828 9090 44884 9100
rect 44604 8866 44660 8876
rect 44716 8930 44772 8942
rect 44716 8878 44718 8930
rect 44770 8878 44772 8930
rect 43932 8820 43988 8830
rect 43932 8726 43988 8764
rect 44268 8818 44324 8830
rect 44268 8766 44270 8818
rect 44322 8766 44324 8818
rect 42812 7308 43092 7364
rect 43708 8484 43764 8494
rect 42476 7252 42532 7262
rect 42532 7196 42644 7252
rect 42476 7186 42532 7196
rect 42588 6690 42644 7196
rect 42588 6638 42590 6690
rect 42642 6638 42644 6690
rect 42588 6626 42644 6638
rect 42812 6690 42868 7308
rect 42812 6638 42814 6690
rect 42866 6638 42868 6690
rect 42812 6468 42868 6638
rect 43484 6692 43540 6702
rect 43708 6692 43764 8428
rect 43932 7474 43988 7486
rect 43932 7422 43934 7474
rect 43986 7422 43988 7474
rect 43932 7364 43988 7422
rect 44268 7476 44324 8766
rect 44268 7410 44324 7420
rect 44604 7476 44660 7486
rect 44716 7476 44772 8878
rect 44940 8932 44996 8942
rect 44940 8482 44996 8876
rect 44940 8430 44942 8482
rect 44994 8430 44996 8482
rect 44940 8418 44996 8430
rect 45276 8484 45332 9212
rect 45276 8370 45332 8428
rect 45276 8318 45278 8370
rect 45330 8318 45332 8370
rect 45276 8306 45332 8318
rect 45500 8372 45556 10334
rect 45724 9940 45780 11452
rect 45836 14588 46116 14644
rect 46396 14644 46452 14654
rect 46396 14642 46676 14644
rect 46396 14590 46398 14642
rect 46450 14590 46676 14642
rect 46396 14588 46676 14590
rect 45836 10836 45892 14588
rect 46396 14578 46452 14588
rect 46284 14530 46340 14542
rect 46284 14478 46286 14530
rect 46338 14478 46340 14530
rect 45948 14420 46004 14430
rect 46284 14420 46340 14478
rect 45948 14418 46340 14420
rect 45948 14366 45950 14418
rect 46002 14366 46340 14418
rect 45948 14364 46340 14366
rect 45948 14354 46004 14364
rect 46508 14308 46564 14318
rect 46508 14214 46564 14252
rect 46284 14196 46340 14206
rect 46060 13860 46116 13870
rect 46060 13766 46116 13804
rect 46172 12292 46228 12302
rect 46172 12198 46228 12236
rect 45948 10836 46004 10846
rect 45836 10834 46004 10836
rect 45836 10782 45950 10834
rect 46002 10782 46004 10834
rect 45836 10780 46004 10782
rect 45836 10388 45892 10780
rect 45948 10770 46004 10780
rect 45836 10322 45892 10332
rect 46284 10500 46340 14140
rect 46620 12964 46676 14588
rect 46732 14420 46788 14430
rect 46732 14326 46788 14364
rect 46844 13076 46900 15092
rect 47180 14530 47236 15092
rect 47180 14478 47182 14530
rect 47234 14478 47236 14530
rect 47180 13860 47236 14478
rect 47404 14530 47460 17276
rect 47516 16100 47572 16110
rect 47740 16100 47796 18396
rect 48972 18452 49028 18462
rect 48972 17778 49028 18396
rect 49196 18338 49252 21084
rect 49420 20914 49476 21644
rect 49756 21588 49812 21598
rect 49420 20862 49422 20914
rect 49474 20862 49476 20914
rect 49420 20580 49476 20862
rect 49420 20514 49476 20524
rect 49644 21586 49812 21588
rect 49644 21534 49758 21586
rect 49810 21534 49812 21586
rect 49644 21532 49812 21534
rect 49644 20802 49700 21532
rect 49756 21522 49812 21532
rect 49980 21026 50036 21868
rect 49980 20974 49982 21026
rect 50034 20974 50036 21026
rect 49980 20962 50036 20974
rect 50540 21812 50596 21822
rect 50540 20916 50596 21756
rect 50876 21586 50932 22428
rect 50876 21534 50878 21586
rect 50930 21534 50932 21586
rect 50876 21522 50932 21534
rect 50540 20822 50596 20860
rect 49644 20750 49646 20802
rect 49698 20750 49700 20802
rect 49644 20692 49700 20750
rect 50988 20802 51044 22652
rect 52948 22652 53172 22708
rect 52892 22642 52948 22652
rect 53116 22372 53172 22652
rect 53116 21586 53172 22316
rect 53116 21534 53118 21586
rect 53170 21534 53172 21586
rect 53116 21522 53172 21534
rect 53228 22260 53284 23100
rect 53452 22260 53508 23886
rect 53564 23156 53620 24220
rect 53676 24162 53732 26012
rect 55020 25508 55076 26350
rect 57932 26292 57988 26302
rect 57932 25730 57988 26236
rect 57932 25678 57934 25730
rect 57986 25678 57988 25730
rect 57932 25666 57988 25678
rect 55580 25508 55636 25518
rect 55020 25506 55636 25508
rect 55020 25454 55582 25506
rect 55634 25454 55636 25506
rect 55020 25452 55636 25454
rect 55580 25442 55636 25452
rect 57932 24948 57988 24958
rect 53900 24724 53956 24734
rect 53900 24722 54516 24724
rect 53900 24670 53902 24722
rect 53954 24670 54516 24722
rect 53900 24668 54516 24670
rect 53900 24658 53956 24668
rect 53676 24110 53678 24162
rect 53730 24110 53732 24162
rect 53676 24098 53732 24110
rect 54460 23826 54516 24668
rect 55356 24498 55412 24510
rect 55356 24446 55358 24498
rect 55410 24446 55412 24498
rect 55356 24276 55412 24446
rect 55356 24210 55412 24220
rect 57932 24162 57988 24892
rect 57932 24110 57934 24162
rect 57986 24110 57988 24162
rect 57932 24098 57988 24110
rect 54684 23940 54740 23950
rect 54460 23774 54462 23826
rect 54514 23774 54516 23826
rect 54460 23762 54516 23774
rect 54572 23938 54740 23940
rect 54572 23886 54686 23938
rect 54738 23886 54740 23938
rect 54572 23884 54740 23886
rect 54460 23268 54516 23278
rect 54572 23268 54628 23884
rect 54684 23874 54740 23884
rect 55580 23940 55636 23950
rect 55580 23846 55636 23884
rect 54460 23266 54628 23268
rect 54460 23214 54462 23266
rect 54514 23214 54628 23266
rect 54460 23212 54628 23214
rect 54460 23202 54516 23212
rect 53788 23156 53844 23166
rect 53564 23154 53844 23156
rect 53564 23102 53790 23154
rect 53842 23102 53844 23154
rect 53564 23100 53844 23102
rect 53788 23090 53844 23100
rect 54012 23042 54068 23054
rect 54012 22990 54014 23042
rect 54066 22990 54068 23042
rect 54012 22596 54068 22990
rect 53788 22540 54068 22596
rect 53788 22482 53844 22540
rect 54348 22484 54404 22494
rect 53788 22430 53790 22482
rect 53842 22430 53844 22482
rect 53788 22418 53844 22430
rect 53900 22482 54404 22484
rect 53900 22430 54350 22482
rect 54402 22430 54404 22482
rect 53900 22428 54404 22430
rect 53900 22370 53956 22428
rect 54348 22418 54404 22428
rect 53900 22318 53902 22370
rect 53954 22318 53956 22370
rect 53900 22306 53956 22318
rect 54460 22372 54516 22382
rect 53564 22260 53620 22270
rect 53452 22258 53620 22260
rect 53452 22206 53566 22258
rect 53618 22206 53620 22258
rect 53452 22204 53620 22206
rect 51660 21474 51716 21486
rect 51660 21422 51662 21474
rect 51714 21422 51716 21474
rect 51548 21364 51604 21374
rect 50988 20750 50990 20802
rect 51042 20750 51044 20802
rect 50988 20738 51044 20750
rect 51212 20916 51268 20926
rect 51212 20802 51268 20860
rect 51212 20750 51214 20802
rect 51266 20750 51268 20802
rect 51212 20738 51268 20750
rect 50316 20692 50372 20702
rect 49644 20690 50372 20692
rect 49644 20638 50318 20690
rect 50370 20638 50372 20690
rect 49644 20636 50372 20638
rect 49644 20132 49700 20636
rect 50316 20626 50372 20636
rect 50540 20580 50596 20618
rect 50540 20514 50596 20524
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 49644 20066 49700 20076
rect 50764 19236 50820 19246
rect 51324 19236 51380 19246
rect 50428 19234 51380 19236
rect 50428 19182 50766 19234
rect 50818 19182 51326 19234
rect 51378 19182 51380 19234
rect 50428 19180 51380 19182
rect 49196 18286 49198 18338
rect 49250 18286 49252 18338
rect 49196 17890 49252 18286
rect 49196 17838 49198 17890
rect 49250 17838 49252 17890
rect 49196 17826 49252 17838
rect 49532 18452 49588 18462
rect 49532 17890 49588 18396
rect 49868 18452 49924 18462
rect 50428 18452 50484 19180
rect 50764 19170 50820 19180
rect 51324 19170 51380 19180
rect 51548 19234 51604 21308
rect 51548 19182 51550 19234
rect 51602 19182 51604 19234
rect 50540 19012 50596 19050
rect 50540 18946 50596 18956
rect 50876 19010 50932 19022
rect 50876 18958 50878 19010
rect 50930 18958 50932 19010
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50876 18676 50932 18958
rect 49868 18450 50484 18452
rect 49868 18398 49870 18450
rect 49922 18398 50484 18450
rect 49868 18396 50484 18398
rect 49868 18386 49924 18396
rect 49532 17838 49534 17890
rect 49586 17838 49588 17890
rect 49532 17826 49588 17838
rect 48972 17726 48974 17778
rect 49026 17726 49028 17778
rect 48972 17714 49028 17726
rect 50428 17666 50484 18396
rect 50764 18620 50932 18676
rect 50988 19012 51044 19022
rect 51548 19012 51604 19182
rect 50988 19010 51604 19012
rect 50988 18958 50990 19010
rect 51042 18958 51604 19010
rect 50988 18956 51604 18958
rect 50764 18338 50820 18620
rect 50764 18286 50766 18338
rect 50818 18286 50820 18338
rect 50764 18274 50820 18286
rect 50428 17614 50430 17666
rect 50482 17614 50484 17666
rect 50428 17602 50484 17614
rect 50988 17666 51044 18956
rect 51100 18452 51156 18462
rect 51100 18358 51156 18396
rect 51660 18452 51716 21422
rect 53228 21476 53284 22204
rect 53340 21476 53396 21486
rect 53228 21474 53396 21476
rect 53228 21422 53342 21474
rect 53394 21422 53396 21474
rect 53228 21420 53396 21422
rect 51772 20916 51828 20926
rect 51772 20822 51828 20860
rect 53340 20916 53396 21420
rect 53564 21476 53620 22204
rect 54236 22260 54292 22270
rect 54236 22166 54292 22204
rect 54460 22258 54516 22316
rect 54460 22206 54462 22258
rect 54514 22206 54516 22258
rect 54460 22194 54516 22206
rect 53564 21410 53620 21420
rect 54012 21700 54068 21710
rect 54572 21700 54628 21710
rect 54012 21698 54628 21700
rect 54012 21646 54014 21698
rect 54066 21646 54574 21698
rect 54626 21646 54628 21698
rect 54012 21644 54628 21646
rect 53340 20850 53396 20860
rect 54012 20802 54068 21644
rect 54572 21634 54628 21644
rect 54460 21476 54516 21486
rect 54460 21382 54516 21420
rect 54348 21362 54404 21374
rect 54348 21310 54350 21362
rect 54402 21310 54404 21362
rect 54012 20750 54014 20802
rect 54066 20750 54068 20802
rect 54012 20738 54068 20750
rect 54236 20804 54292 20814
rect 54348 20804 54404 21310
rect 57932 20916 57988 20926
rect 57932 20822 57988 20860
rect 55580 20804 55636 20814
rect 54236 20802 54404 20804
rect 54236 20750 54238 20802
rect 54290 20750 54404 20802
rect 54236 20748 54404 20750
rect 55132 20802 55636 20804
rect 55132 20750 55582 20802
rect 55634 20750 55636 20802
rect 55132 20748 55636 20750
rect 51884 19346 51940 19358
rect 51884 19294 51886 19346
rect 51938 19294 51940 19346
rect 51884 19236 51940 19294
rect 51884 19170 51940 19180
rect 53228 19236 53284 19246
rect 53284 19180 53508 19236
rect 53228 19142 53284 19180
rect 52892 19122 52948 19134
rect 52892 19070 52894 19122
rect 52946 19070 52948 19122
rect 52892 19012 52948 19070
rect 51996 18564 52052 18574
rect 51996 18562 52164 18564
rect 51996 18510 51998 18562
rect 52050 18510 52164 18562
rect 51996 18508 52164 18510
rect 51996 18498 52052 18508
rect 51660 18386 51716 18396
rect 50988 17614 50990 17666
rect 51042 17614 51044 17666
rect 50988 17602 51044 17614
rect 51548 18338 51604 18350
rect 51548 18286 51550 18338
rect 51602 18286 51604 18338
rect 51100 17554 51156 17566
rect 51100 17502 51102 17554
rect 51154 17502 51156 17554
rect 47572 16044 47796 16100
rect 47964 17444 48020 17454
rect 47964 17108 48020 17388
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 47964 16098 48020 17052
rect 47964 16046 47966 16098
rect 48018 16046 48020 16098
rect 47516 16006 47572 16044
rect 47964 16034 48020 16046
rect 48188 16660 48244 16670
rect 48188 16098 48244 16604
rect 49532 16212 49588 16222
rect 49532 16118 49588 16156
rect 50092 16212 50148 16222
rect 48188 16046 48190 16098
rect 48242 16046 48244 16098
rect 48188 16034 48244 16046
rect 48076 15876 48132 15886
rect 48076 15782 48132 15820
rect 49084 15876 49140 15886
rect 49084 15314 49140 15820
rect 49644 15876 49700 15886
rect 49644 15782 49700 15820
rect 49084 15262 49086 15314
rect 49138 15262 49140 15314
rect 48860 15202 48916 15214
rect 48860 15150 48862 15202
rect 48914 15150 48916 15202
rect 48860 15148 48916 15150
rect 47404 14478 47406 14530
rect 47458 14478 47460 14530
rect 47404 14466 47460 14478
rect 48748 15092 48916 15148
rect 48748 14530 48804 15092
rect 48860 15026 48916 15036
rect 49084 15204 49140 15262
rect 49420 15316 49476 15326
rect 49420 15222 49476 15260
rect 49084 14642 49140 15148
rect 49756 15202 49812 15214
rect 49756 15150 49758 15202
rect 49810 15150 49812 15202
rect 49756 15092 49812 15150
rect 49980 15204 50036 15242
rect 49980 15138 50036 15148
rect 49756 15026 49812 15036
rect 49084 14590 49086 14642
rect 49138 14590 49140 14642
rect 49084 14578 49140 14590
rect 48748 14478 48750 14530
rect 48802 14478 48804 14530
rect 47964 14420 48020 14430
rect 47964 14418 48356 14420
rect 47964 14366 47966 14418
rect 48018 14366 48356 14418
rect 47964 14364 48356 14366
rect 47964 14354 48020 14364
rect 47180 13794 47236 13804
rect 46956 13076 47012 13086
rect 46844 13074 47572 13076
rect 46844 13022 46958 13074
rect 47010 13022 47572 13074
rect 46844 13020 47572 13022
rect 46956 13010 47012 13020
rect 46620 12962 46788 12964
rect 46620 12910 46622 12962
rect 46674 12910 46788 12962
rect 46620 12908 46788 12910
rect 46620 12898 46676 12908
rect 46396 11508 46452 11518
rect 46396 11414 46452 11452
rect 46732 11508 46788 12908
rect 47404 12628 47460 12638
rect 46956 12178 47012 12190
rect 46956 12126 46958 12178
rect 47010 12126 47012 12178
rect 46732 11506 46900 11508
rect 46732 11454 46734 11506
rect 46786 11454 46900 11506
rect 46732 11452 46900 11454
rect 46732 11442 46788 11452
rect 46732 10724 46788 10734
rect 46732 10612 46788 10668
rect 46620 10610 46788 10612
rect 46620 10558 46734 10610
rect 46786 10558 46788 10610
rect 46620 10556 46788 10558
rect 46396 10500 46452 10510
rect 46284 10498 46452 10500
rect 46284 10446 46398 10498
rect 46450 10446 46452 10498
rect 46284 10444 46452 10446
rect 45836 9940 45892 9950
rect 45724 9938 45892 9940
rect 45724 9886 45838 9938
rect 45890 9886 45892 9938
rect 45724 9884 45892 9886
rect 45836 9874 45892 9884
rect 45612 9268 45668 9278
rect 45612 9174 45668 9212
rect 46284 9268 46340 10444
rect 46396 10434 46452 10444
rect 46620 9828 46676 10556
rect 46732 10546 46788 10556
rect 46844 10050 46900 11452
rect 46956 11396 47012 12126
rect 47404 12068 47460 12572
rect 47180 12066 47460 12068
rect 47180 12014 47406 12066
rect 47458 12014 47460 12066
rect 47180 12012 47460 12014
rect 47180 11618 47236 12012
rect 47404 12002 47460 12012
rect 47516 12178 47572 13020
rect 47516 12126 47518 12178
rect 47570 12126 47572 12178
rect 47180 11566 47182 11618
rect 47234 11566 47236 11618
rect 47180 11554 47236 11566
rect 47516 11844 47572 12126
rect 48188 12290 48244 12302
rect 48188 12238 48190 12290
rect 48242 12238 48244 12290
rect 48188 12180 48244 12238
rect 48188 12114 48244 12124
rect 46956 11302 47012 11340
rect 47292 10612 47348 10622
rect 46844 9998 46846 10050
rect 46898 9998 46900 10050
rect 46844 9986 46900 9998
rect 47068 10556 47292 10612
rect 47068 10050 47124 10556
rect 47292 10546 47348 10556
rect 47516 10610 47572 11788
rect 48300 11620 48356 14364
rect 48748 12404 48804 14478
rect 50092 14530 50148 16156
rect 50988 16212 51044 16222
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50988 15540 51044 16156
rect 51100 16100 51156 17502
rect 51548 16884 51604 18286
rect 51548 16818 51604 16828
rect 52108 17108 52164 18508
rect 52556 18450 52612 18462
rect 52556 18398 52558 18450
rect 52610 18398 52612 18450
rect 52556 17778 52612 18398
rect 52556 17726 52558 17778
rect 52610 17726 52612 17778
rect 52556 17714 52612 17726
rect 52668 18452 52724 18462
rect 52668 17666 52724 18396
rect 52668 17614 52670 17666
rect 52722 17614 52724 17666
rect 52668 17602 52724 17614
rect 52892 17554 52948 18956
rect 52892 17502 52894 17554
rect 52946 17502 52948 17554
rect 52892 17490 52948 17502
rect 53228 18564 53284 18574
rect 52108 16322 52164 17052
rect 53228 17106 53284 18508
rect 53452 17554 53508 19180
rect 53564 19234 53620 19246
rect 53564 19182 53566 19234
rect 53618 19182 53620 19234
rect 53564 18452 53620 19182
rect 53676 19010 53732 19022
rect 53676 18958 53678 19010
rect 53730 18958 53732 19010
rect 53676 18452 53732 18958
rect 54236 18562 54292 20748
rect 54460 20692 54516 20702
rect 54796 20692 54852 20702
rect 54460 20690 54852 20692
rect 54460 20638 54462 20690
rect 54514 20638 54798 20690
rect 54850 20638 54852 20690
rect 54460 20636 54852 20638
rect 54460 20626 54516 20636
rect 54796 20626 54852 20636
rect 55132 20690 55188 20748
rect 55580 20738 55636 20748
rect 55132 20638 55134 20690
rect 55186 20638 55188 20690
rect 55132 20626 55188 20638
rect 54236 18510 54238 18562
rect 54290 18510 54292 18562
rect 54236 18498 54292 18510
rect 55132 18564 55188 18574
rect 55132 18470 55188 18508
rect 53788 18452 53844 18462
rect 53676 18450 53844 18452
rect 53676 18398 53790 18450
rect 53842 18398 53844 18450
rect 53676 18396 53844 18398
rect 53564 18386 53620 18396
rect 53788 18386 53844 18396
rect 55692 18450 55748 18462
rect 55692 18398 55694 18450
rect 55746 18398 55748 18450
rect 53452 17502 53454 17554
rect 53506 17502 53508 17554
rect 53452 17490 53508 17502
rect 54348 17778 54404 17790
rect 54348 17726 54350 17778
rect 54402 17726 54404 17778
rect 53228 17054 53230 17106
rect 53282 17054 53284 17106
rect 53228 17042 53284 17054
rect 54348 17106 54404 17726
rect 54572 17666 54628 17678
rect 55580 17668 55636 17678
rect 54572 17614 54574 17666
rect 54626 17614 54628 17666
rect 54348 17054 54350 17106
rect 54402 17054 54404 17106
rect 54348 17042 54404 17054
rect 54460 17108 54516 17118
rect 54460 17014 54516 17052
rect 53340 16884 53396 16894
rect 53340 16770 53396 16828
rect 53564 16884 53620 16894
rect 54572 16884 54628 17614
rect 55244 17666 55636 17668
rect 55244 17614 55582 17666
rect 55634 17614 55636 17666
rect 55244 17612 55636 17614
rect 55132 17556 55188 17566
rect 53564 16882 53732 16884
rect 53564 16830 53566 16882
rect 53618 16830 53732 16882
rect 53564 16828 53732 16830
rect 53564 16818 53620 16828
rect 53340 16718 53342 16770
rect 53394 16718 53396 16770
rect 53340 16706 53396 16718
rect 52108 16270 52110 16322
rect 52162 16270 52164 16322
rect 52108 16258 52164 16270
rect 52780 16660 52836 16670
rect 51772 16212 51828 16222
rect 51772 16118 51828 16156
rect 51548 16100 51604 16110
rect 51100 16044 51548 16100
rect 51548 16006 51604 16044
rect 51212 15876 51268 15886
rect 51100 15540 51156 15550
rect 50988 15538 51156 15540
rect 50988 15486 51102 15538
rect 51154 15486 51156 15538
rect 50988 15484 51156 15486
rect 51100 15474 51156 15484
rect 51212 15538 51268 15820
rect 51212 15486 51214 15538
rect 51266 15486 51268 15538
rect 51212 15474 51268 15486
rect 52780 15538 52836 16604
rect 53004 16212 53060 16222
rect 53004 16118 53060 16156
rect 53676 16210 53732 16828
rect 54572 16818 54628 16828
rect 55020 17554 55188 17556
rect 55020 17502 55134 17554
rect 55186 17502 55188 17554
rect 55020 17500 55188 17502
rect 55020 16882 55076 17500
rect 55132 17490 55188 17500
rect 55244 17106 55300 17612
rect 55580 17602 55636 17612
rect 55244 17054 55246 17106
rect 55298 17054 55300 17106
rect 55244 17042 55300 17054
rect 55020 16830 55022 16882
rect 55074 16830 55076 16882
rect 55020 16818 55076 16830
rect 54236 16660 54292 16670
rect 54236 16566 54292 16604
rect 53676 16158 53678 16210
rect 53730 16158 53732 16210
rect 52892 16100 52948 16110
rect 52892 16006 52948 16044
rect 52780 15486 52782 15538
rect 52834 15486 52836 15538
rect 52780 15474 52836 15486
rect 52668 15428 52724 15438
rect 52668 15334 52724 15372
rect 53564 15428 53620 15438
rect 53676 15428 53732 16158
rect 53620 15372 53732 15428
rect 50540 15316 50596 15326
rect 50316 15314 50596 15316
rect 50316 15262 50542 15314
rect 50594 15262 50596 15314
rect 50316 15260 50596 15262
rect 50316 15090 50372 15260
rect 50540 15250 50596 15260
rect 50988 15316 51044 15326
rect 50988 15222 51044 15260
rect 53564 15314 53620 15372
rect 53564 15262 53566 15314
rect 53618 15262 53620 15314
rect 53564 15250 53620 15262
rect 52892 15202 52948 15214
rect 52892 15150 52894 15202
rect 52946 15150 52948 15202
rect 52892 15148 52948 15150
rect 53340 15202 53396 15214
rect 53340 15150 53342 15202
rect 53394 15150 53396 15202
rect 53340 15148 53396 15150
rect 52892 15092 53396 15148
rect 54236 15202 54292 15214
rect 54236 15150 54238 15202
rect 54290 15150 54292 15202
rect 50316 15038 50318 15090
rect 50370 15038 50372 15090
rect 50316 15026 50372 15038
rect 50092 14478 50094 14530
rect 50146 14478 50148 14530
rect 50092 14466 50148 14478
rect 50876 14420 50932 14430
rect 50876 14326 50932 14364
rect 51660 14420 51716 14430
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 51660 13076 51716 14364
rect 52220 14420 52276 14430
rect 51324 12964 51380 12974
rect 51324 12870 51380 12908
rect 51660 12962 51716 13020
rect 51660 12910 51662 12962
rect 51714 12910 51716 12962
rect 51660 12898 51716 12910
rect 51772 13858 51828 13870
rect 51772 13806 51774 13858
rect 51826 13806 51828 13858
rect 51772 12962 51828 13806
rect 52220 13858 52276 14364
rect 52220 13806 52222 13858
rect 52274 13806 52276 13858
rect 52220 13794 52276 13806
rect 51996 13746 52052 13758
rect 51996 13694 51998 13746
rect 52050 13694 52052 13746
rect 51772 12910 51774 12962
rect 51826 12910 51828 12962
rect 49756 12852 49812 12862
rect 49756 12758 49812 12796
rect 50988 12850 51044 12862
rect 50988 12798 50990 12850
rect 51042 12798 51044 12850
rect 48748 12338 48804 12348
rect 49420 12738 49476 12750
rect 49420 12686 49422 12738
rect 49474 12686 49476 12738
rect 48972 12292 49028 12302
rect 48860 12180 48916 12190
rect 48860 12086 48916 12124
rect 48076 11618 48356 11620
rect 48076 11566 48302 11618
rect 48354 11566 48356 11618
rect 48076 11564 48356 11566
rect 47628 11396 47684 11406
rect 47628 11302 47684 11340
rect 47964 11394 48020 11406
rect 47964 11342 47966 11394
rect 48018 11342 48020 11394
rect 47516 10558 47518 10610
rect 47570 10558 47572 10610
rect 47516 10546 47572 10558
rect 47852 11282 47908 11294
rect 47852 11230 47854 11282
rect 47906 11230 47908 11282
rect 47068 9998 47070 10050
rect 47122 9998 47124 10050
rect 47068 9986 47124 9998
rect 46620 9734 46676 9772
rect 47852 9826 47908 11230
rect 47964 10724 48020 11342
rect 47964 10658 48020 10668
rect 48076 10612 48132 11564
rect 48300 11554 48356 11564
rect 48412 11844 48468 11854
rect 48188 11396 48244 11406
rect 48412 11396 48468 11788
rect 48188 11394 48468 11396
rect 48188 11342 48190 11394
rect 48242 11342 48468 11394
rect 48188 11340 48468 11342
rect 48972 11396 49028 12236
rect 49084 12290 49140 12302
rect 49084 12238 49086 12290
rect 49138 12238 49140 12290
rect 49084 11844 49140 12238
rect 49308 12292 49364 12302
rect 49308 12198 49364 12236
rect 49420 11844 49476 12686
rect 50988 12740 51044 12798
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50204 12404 50260 12414
rect 49980 12292 50036 12302
rect 49980 12198 50036 12236
rect 49084 11788 49476 11844
rect 49532 12180 49588 12190
rect 49084 11396 49140 11406
rect 48972 11394 49140 11396
rect 48972 11342 49086 11394
rect 49138 11342 49140 11394
rect 48972 11340 49140 11342
rect 48188 11330 48244 11340
rect 49084 11330 49140 11340
rect 49308 11396 49364 11788
rect 49308 11302 49364 11340
rect 49420 11396 49476 11406
rect 49532 11396 49588 12124
rect 50204 12178 50260 12348
rect 50204 12126 50206 12178
rect 50258 12126 50260 12178
rect 50204 12114 50260 12126
rect 50428 12402 50484 12414
rect 50428 12350 50430 12402
rect 50482 12350 50484 12402
rect 49420 11394 49588 11396
rect 49420 11342 49422 11394
rect 49474 11342 49588 11394
rect 49420 11340 49588 11342
rect 49420 11330 49476 11340
rect 49868 11172 49924 11182
rect 49868 11170 50148 11172
rect 49868 11118 49870 11170
rect 49922 11118 50148 11170
rect 49868 11116 50148 11118
rect 49868 11106 49924 11116
rect 50092 10834 50148 11116
rect 50092 10782 50094 10834
rect 50146 10782 50148 10834
rect 48188 10724 48244 10734
rect 48188 10722 48468 10724
rect 48188 10670 48190 10722
rect 48242 10670 48468 10722
rect 48188 10668 48468 10670
rect 48188 10658 48244 10668
rect 48076 10518 48132 10556
rect 47852 9774 47854 9826
rect 47906 9774 47908 9826
rect 47852 9762 47908 9774
rect 48412 9826 48468 10668
rect 48636 10612 48692 10622
rect 48636 9938 48692 10556
rect 49644 10612 49700 10622
rect 49644 10518 49700 10556
rect 50092 10388 50148 10782
rect 50316 10836 50372 10846
rect 50428 10836 50484 12350
rect 50988 12292 51044 12684
rect 50988 12226 51044 12236
rect 51100 12852 51156 12862
rect 51100 12290 51156 12796
rect 51772 12852 51828 12910
rect 51772 12786 51828 12796
rect 51884 13634 51940 13646
rect 51884 13582 51886 13634
rect 51938 13582 51940 13634
rect 51884 12404 51940 13582
rect 51996 12964 52052 13694
rect 52780 13076 52836 13086
rect 52780 12982 52836 13020
rect 53004 12964 53060 12974
rect 51996 12908 52164 12964
rect 52108 12850 52164 12908
rect 53004 12870 53060 12908
rect 52108 12798 52110 12850
rect 52162 12798 52164 12850
rect 51996 12738 52052 12750
rect 51996 12686 51998 12738
rect 52050 12686 52052 12738
rect 51996 12516 52052 12686
rect 52108 12740 52164 12798
rect 52108 12674 52164 12684
rect 51996 12460 52388 12516
rect 51884 12310 51940 12348
rect 52332 12402 52388 12460
rect 52332 12350 52334 12402
rect 52386 12350 52388 12402
rect 51100 12238 51102 12290
rect 51154 12238 51156 12290
rect 51100 12226 51156 12238
rect 50764 12180 50820 12190
rect 50764 12086 50820 12124
rect 52108 12178 52164 12190
rect 52108 12126 52110 12178
rect 52162 12126 52164 12178
rect 52108 11732 52164 12126
rect 52332 12180 52388 12350
rect 52668 12404 52724 12414
rect 52668 12290 52724 12348
rect 52668 12238 52670 12290
rect 52722 12238 52724 12290
rect 52668 12226 52724 12238
rect 53004 12292 53060 12302
rect 53116 12292 53172 15092
rect 54236 14530 54292 15150
rect 54236 14478 54238 14530
rect 54290 14478 54292 14530
rect 54236 14466 54292 14478
rect 54572 14532 54628 14542
rect 54572 14418 54628 14476
rect 55580 14532 55636 14542
rect 55580 14438 55636 14476
rect 54572 14366 54574 14418
rect 54626 14366 54628 14418
rect 54572 14354 54628 14366
rect 53004 12290 53172 12292
rect 53004 12238 53006 12290
rect 53058 12238 53172 12290
rect 53004 12236 53172 12238
rect 53676 12850 53732 12862
rect 53676 12798 53678 12850
rect 53730 12798 53732 12850
rect 53004 12226 53060 12236
rect 52332 12114 52388 12124
rect 52780 12178 52836 12190
rect 52780 12126 52782 12178
rect 52834 12126 52836 12178
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50316 10834 50484 10836
rect 50316 10782 50318 10834
rect 50370 10782 50484 10834
rect 50316 10780 50484 10782
rect 50316 10770 50372 10780
rect 50428 10612 50484 10780
rect 51996 10836 52052 10846
rect 52108 10836 52164 11676
rect 52220 12066 52276 12078
rect 52220 12014 52222 12066
rect 52274 12014 52276 12066
rect 52220 11396 52276 12014
rect 52780 11732 52836 12126
rect 53452 12180 53508 12190
rect 53676 12180 53732 12798
rect 53900 12180 53956 12190
rect 53676 12124 53900 12180
rect 53452 12086 53508 12124
rect 52780 11666 52836 11676
rect 53228 11954 53284 11966
rect 53228 11902 53230 11954
rect 53282 11902 53284 11954
rect 53004 11508 53060 11518
rect 52220 11330 52276 11340
rect 52668 11506 53060 11508
rect 52668 11454 53006 11506
rect 53058 11454 53060 11506
rect 52668 11452 53060 11454
rect 51996 10834 52164 10836
rect 51996 10782 51998 10834
rect 52050 10782 52164 10834
rect 51996 10780 52164 10782
rect 51996 10770 52052 10780
rect 51100 10612 51156 10622
rect 50484 10556 50708 10612
rect 50428 10546 50484 10556
rect 50092 10322 50148 10332
rect 50204 10498 50260 10510
rect 50204 10446 50206 10498
rect 50258 10446 50260 10498
rect 48636 9886 48638 9938
rect 48690 9886 48692 9938
rect 48636 9874 48692 9886
rect 48412 9774 48414 9826
rect 48466 9774 48468 9826
rect 47516 9604 47572 9614
rect 47516 9602 47908 9604
rect 47516 9550 47518 9602
rect 47570 9550 47908 9602
rect 47516 9548 47908 9550
rect 47516 9538 47572 9548
rect 46284 9202 46340 9212
rect 47852 9156 47908 9548
rect 48412 9268 48468 9774
rect 48972 9714 49028 9726
rect 48972 9662 48974 9714
rect 49026 9662 49028 9714
rect 48972 9268 49028 9662
rect 50204 9716 50260 10446
rect 50540 10388 50596 10398
rect 50540 9938 50596 10332
rect 50652 10052 50708 10556
rect 51100 10518 51156 10556
rect 51212 10610 51268 10622
rect 51212 10558 51214 10610
rect 51266 10558 51268 10610
rect 50764 10500 50820 10510
rect 50820 10444 51044 10500
rect 50764 10406 50820 10444
rect 50764 10052 50820 10062
rect 50652 10050 50820 10052
rect 50652 9998 50766 10050
rect 50818 9998 50820 10050
rect 50652 9996 50820 9998
rect 50764 9986 50820 9996
rect 50988 10050 51044 10444
rect 51212 10388 51268 10558
rect 52668 10500 52724 11452
rect 53004 11442 53060 11452
rect 52780 11282 52836 11294
rect 52780 11230 52782 11282
rect 52834 11230 52836 11282
rect 52780 10724 52836 11230
rect 53004 10724 53060 10734
rect 52780 10722 53060 10724
rect 52780 10670 53006 10722
rect 53058 10670 53060 10722
rect 52780 10668 53060 10670
rect 52780 10500 52836 10510
rect 51212 10322 51268 10332
rect 52556 10498 52836 10500
rect 52556 10446 52782 10498
rect 52834 10446 52836 10498
rect 52556 10444 52836 10446
rect 50988 9998 50990 10050
rect 51042 9998 51044 10050
rect 50988 9986 51044 9998
rect 50540 9886 50542 9938
rect 50594 9886 50596 9938
rect 50540 9874 50596 9886
rect 51436 9940 51492 9950
rect 51436 9938 51828 9940
rect 51436 9886 51438 9938
rect 51490 9886 51828 9938
rect 51436 9884 51828 9886
rect 51436 9874 51492 9884
rect 50204 9650 50260 9660
rect 51660 9716 51716 9726
rect 51660 9622 51716 9660
rect 51772 9714 51828 9884
rect 51772 9662 51774 9714
rect 51826 9662 51828 9714
rect 51772 9650 51828 9662
rect 51996 9602 52052 9614
rect 51996 9550 51998 9602
rect 52050 9550 52052 9602
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 48412 9212 48804 9268
rect 48972 9212 49588 9268
rect 45500 8306 45556 8316
rect 47740 8372 47796 8382
rect 45052 8258 45108 8270
rect 45052 8206 45054 8258
rect 45106 8206 45108 8258
rect 45052 7588 45108 8206
rect 47740 8258 47796 8316
rect 47740 8206 47742 8258
rect 47794 8206 47796 8258
rect 45388 8148 45444 8158
rect 45724 8148 45780 8158
rect 45948 8148 46004 8158
rect 45388 8146 45780 8148
rect 45388 8094 45390 8146
rect 45442 8094 45726 8146
rect 45778 8094 45780 8146
rect 45388 8092 45780 8094
rect 45388 8082 45444 8092
rect 45724 8082 45780 8092
rect 45836 8146 46004 8148
rect 45836 8094 45950 8146
rect 46002 8094 46004 8146
rect 45836 8092 46004 8094
rect 45052 7532 45332 7588
rect 44604 7474 45220 7476
rect 44604 7422 44606 7474
rect 44658 7422 45220 7474
rect 44604 7420 45220 7422
rect 44604 7410 44660 7420
rect 43932 7298 43988 7308
rect 45164 6802 45220 7420
rect 45164 6750 45166 6802
rect 45218 6750 45220 6802
rect 45164 6738 45220 6750
rect 45276 7364 45332 7532
rect 45500 7476 45556 7486
rect 45500 7382 45556 7420
rect 43540 6636 43764 6692
rect 45276 6690 45332 7308
rect 45836 6914 45892 8092
rect 45948 8082 46004 8092
rect 46284 8146 46340 8158
rect 46284 8094 46286 8146
rect 46338 8094 46340 8146
rect 46172 8034 46228 8046
rect 46172 7982 46174 8034
rect 46226 7982 46228 8034
rect 45836 6862 45838 6914
rect 45890 6862 45892 6914
rect 45836 6850 45892 6862
rect 46060 7362 46116 7374
rect 46060 7310 46062 7362
rect 46114 7310 46116 7362
rect 45276 6638 45278 6690
rect 45330 6638 45332 6690
rect 43484 6598 43540 6636
rect 45276 6626 45332 6638
rect 42140 5954 42196 5964
rect 42364 6412 42868 6468
rect 42028 5854 42030 5906
rect 42082 5854 42084 5906
rect 42028 5842 42084 5854
rect 42364 5906 42420 6412
rect 46060 6132 46116 7310
rect 46172 7252 46228 7982
rect 46284 7476 46340 8094
rect 46284 7410 46340 7420
rect 46172 7186 46228 7196
rect 47740 6802 47796 8206
rect 47852 8258 47908 9100
rect 47852 8206 47854 8258
rect 47906 8206 47908 8258
rect 47852 8194 47908 8206
rect 47964 8260 48020 8270
rect 48636 8260 48692 9212
rect 48748 9154 48804 9212
rect 48748 9102 48750 9154
rect 48802 9102 48804 9154
rect 48748 9090 48804 9102
rect 48860 9156 48916 9166
rect 48916 9100 49028 9156
rect 48860 9062 48916 9100
rect 47964 8258 48692 8260
rect 47964 8206 47966 8258
rect 48018 8206 48638 8258
rect 48690 8206 48692 8258
rect 47964 8204 48692 8206
rect 47964 8194 48020 8204
rect 48636 8194 48692 8204
rect 48972 8258 49028 9100
rect 49084 9044 49140 9054
rect 49084 9042 49476 9044
rect 49084 8990 49086 9042
rect 49138 8990 49476 9042
rect 49084 8988 49476 8990
rect 49084 8978 49140 8988
rect 48972 8206 48974 8258
rect 49026 8206 49028 8258
rect 48972 8194 49028 8206
rect 49308 8372 49364 8382
rect 49308 8258 49364 8316
rect 49308 8206 49310 8258
rect 49362 8206 49364 8258
rect 49308 8194 49364 8206
rect 48412 8036 48468 8046
rect 48412 7942 48468 7980
rect 48860 8034 48916 8046
rect 48860 7982 48862 8034
rect 48914 7982 48916 8034
rect 48860 7474 48916 7982
rect 48860 7422 48862 7474
rect 48914 7422 48916 7474
rect 48860 7410 48916 7422
rect 48972 8036 49028 8046
rect 48972 7474 49028 7980
rect 48972 7422 48974 7474
rect 49026 7422 49028 7474
rect 48972 7410 49028 7422
rect 49308 7476 49364 7486
rect 49308 7382 49364 7420
rect 47740 6750 47742 6802
rect 47794 6750 47796 6802
rect 47740 6738 47796 6750
rect 47964 7252 48020 7262
rect 46732 6580 46788 6590
rect 46732 6244 46788 6524
rect 47964 6578 48020 7196
rect 49196 7252 49252 7262
rect 49196 7158 49252 7196
rect 49420 6690 49476 8988
rect 49532 8372 49588 9212
rect 51996 9044 52052 9550
rect 51996 8978 52052 8988
rect 49532 8306 49588 8316
rect 51548 8932 51604 8942
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 51548 7698 51604 8876
rect 52556 8932 52612 10444
rect 52780 10434 52836 10444
rect 52668 9044 52724 9054
rect 53004 9044 53060 10668
rect 53228 10724 53284 11902
rect 53788 11732 53844 11742
rect 53788 10834 53844 11676
rect 53900 11506 53956 12124
rect 54572 12180 54628 12190
rect 54572 12086 54628 12124
rect 55244 12180 55300 12190
rect 55580 12180 55636 12190
rect 55244 12178 55636 12180
rect 55244 12126 55246 12178
rect 55298 12126 55582 12178
rect 55634 12126 55636 12178
rect 55244 12124 55636 12126
rect 55244 12114 55300 12124
rect 55580 12114 55636 12124
rect 54348 12068 54404 12078
rect 53900 11454 53902 11506
rect 53954 11454 53956 11506
rect 53900 11442 53956 11454
rect 54012 12066 54404 12068
rect 54012 12014 54350 12066
rect 54402 12014 54404 12066
rect 54012 12012 54404 12014
rect 53788 10782 53790 10834
rect 53842 10782 53844 10834
rect 53788 10770 53844 10782
rect 53564 10724 53620 10734
rect 53228 10722 53620 10724
rect 53228 10670 53566 10722
rect 53618 10670 53620 10722
rect 53228 10668 53620 10670
rect 53116 10500 53172 10510
rect 53228 10500 53284 10668
rect 53564 10658 53620 10668
rect 53116 10498 53284 10500
rect 53116 10446 53118 10498
rect 53170 10446 53284 10498
rect 53116 10444 53284 10446
rect 53900 10500 53956 10510
rect 54012 10500 54068 12012
rect 54348 12002 54404 12012
rect 54348 11844 54404 11854
rect 54348 11618 54404 11788
rect 55692 11844 55748 18398
rect 57932 17778 57988 17790
rect 57932 17726 57934 17778
rect 57986 17726 57988 17778
rect 57932 17556 57988 17726
rect 57932 17490 57988 17500
rect 57932 14868 57988 14878
rect 57932 14754 57988 14812
rect 57932 14702 57934 14754
rect 57986 14702 57988 14754
rect 57932 14690 57988 14702
rect 57932 13074 57988 13086
rect 57932 13022 57934 13074
rect 57986 13022 57988 13074
rect 55916 12962 55972 12974
rect 55916 12910 55918 12962
rect 55970 12910 55972 12962
rect 55916 12402 55972 12910
rect 55916 12350 55918 12402
rect 55970 12350 55972 12402
rect 55916 12338 55972 12350
rect 57932 12180 57988 13022
rect 57932 12114 57988 12124
rect 55692 11778 55748 11788
rect 54348 11566 54350 11618
rect 54402 11566 54404 11618
rect 54348 11554 54404 11566
rect 54236 11396 54292 11406
rect 54236 11302 54292 11340
rect 53900 10498 54068 10500
rect 53900 10446 53902 10498
rect 53954 10446 54068 10498
rect 53900 10444 54068 10446
rect 53116 10434 53172 10444
rect 53900 10434 53956 10444
rect 54012 9154 54068 9166
rect 54012 9102 54014 9154
rect 54066 9102 54068 9154
rect 52724 8988 53060 9044
rect 53340 9044 53396 9054
rect 53676 9044 53732 9054
rect 53340 9042 53732 9044
rect 53340 8990 53342 9042
rect 53394 8990 53678 9042
rect 53730 8990 53732 9042
rect 53340 8988 53732 8990
rect 52668 8950 52724 8988
rect 53340 8978 53396 8988
rect 53676 8978 53732 8988
rect 52556 8838 52612 8876
rect 54012 8260 54068 9102
rect 57932 8372 57988 8382
rect 57932 8278 57988 8316
rect 54012 8194 54068 8204
rect 55580 8260 55636 8270
rect 55580 8166 55636 8204
rect 51548 7646 51550 7698
rect 51602 7646 51604 7698
rect 51548 7634 51604 7646
rect 50652 7586 50708 7598
rect 50652 7534 50654 7586
rect 50706 7534 50708 7586
rect 50540 7474 50596 7486
rect 50540 7422 50542 7474
rect 50594 7422 50596 7474
rect 49420 6638 49422 6690
rect 49474 6638 49476 6690
rect 49420 6626 49476 6638
rect 49868 6804 49924 6814
rect 49868 6690 49924 6748
rect 50540 6804 50596 7422
rect 50540 6710 50596 6748
rect 49868 6638 49870 6690
rect 49922 6638 49924 6690
rect 49868 6626 49924 6638
rect 50652 6692 50708 7534
rect 51436 7476 51492 7486
rect 51436 7382 51492 7420
rect 50652 6598 50708 6636
rect 47964 6526 47966 6578
rect 48018 6526 48020 6578
rect 47964 6514 48020 6526
rect 51324 6580 51380 6590
rect 51660 6580 51716 6590
rect 51324 6578 51716 6580
rect 51324 6526 51326 6578
rect 51378 6526 51662 6578
rect 51714 6526 51716 6578
rect 51324 6524 51716 6526
rect 51324 6514 51380 6524
rect 51660 6514 51716 6524
rect 51996 6468 52052 6478
rect 51996 6466 52164 6468
rect 51996 6414 51998 6466
rect 52050 6414 52164 6466
rect 51996 6412 52164 6414
rect 51996 6402 52052 6412
rect 47964 6356 48020 6366
rect 46732 6188 47348 6244
rect 46060 6076 46564 6132
rect 46508 6020 46564 6076
rect 46508 5926 46564 5964
rect 46732 6130 46788 6188
rect 46732 6078 46734 6130
rect 46786 6078 46788 6130
rect 42364 5854 42366 5906
rect 42418 5854 42420 5906
rect 42364 5842 42420 5854
rect 42588 5906 42644 5918
rect 42588 5854 42590 5906
rect 42642 5854 42644 5906
rect 42588 5124 42644 5854
rect 46620 5794 46676 5806
rect 46620 5742 46622 5794
rect 46674 5742 46676 5794
rect 42588 5058 42644 5068
rect 42812 5236 42868 5246
rect 42812 5122 42868 5180
rect 45388 5236 45444 5246
rect 42812 5070 42814 5122
rect 42866 5070 42868 5122
rect 42812 5058 42868 5070
rect 43372 5124 43428 5134
rect 43372 5030 43428 5068
rect 43484 5124 43540 5134
rect 43820 5124 43876 5134
rect 43484 5122 43876 5124
rect 43484 5070 43486 5122
rect 43538 5070 43822 5122
rect 43874 5070 43876 5122
rect 43484 5068 43876 5070
rect 43484 5058 43540 5068
rect 43820 5058 43876 5068
rect 45164 5124 45220 5134
rect 45164 5030 45220 5068
rect 41244 4918 41300 4956
rect 45388 5010 45444 5180
rect 45388 4958 45390 5010
rect 45442 4958 45444 5010
rect 45388 4946 45444 4958
rect 45500 5234 45556 5246
rect 45500 5182 45502 5234
rect 45554 5182 45556 5234
rect 45500 5012 45556 5182
rect 46172 5236 46228 5246
rect 46228 5180 46340 5236
rect 46172 5170 46228 5180
rect 46172 5012 46228 5022
rect 45500 5010 46228 5012
rect 45500 4958 46174 5010
rect 46226 4958 46228 5010
rect 45500 4956 46228 4958
rect 46172 4946 46228 4956
rect 44156 4898 44212 4910
rect 44156 4846 44158 4898
rect 44210 4846 44212 4898
rect 40908 4450 40964 4462
rect 40908 4398 40910 4450
rect 40962 4398 40964 4450
rect 40348 4340 40404 4350
rect 40348 4246 40404 4284
rect 39900 4228 39956 4238
rect 39788 4226 39956 4228
rect 39788 4174 39902 4226
rect 39954 4174 39956 4226
rect 39788 4172 39956 4174
rect 39900 4162 39956 4172
rect 40908 3554 40964 4398
rect 41132 4340 41188 4350
rect 41132 4246 41188 4284
rect 40908 3502 40910 3554
rect 40962 3502 40964 3554
rect 40908 3490 40964 3502
rect 44156 3554 44212 4846
rect 46284 4450 46340 5180
rect 46284 4398 46286 4450
rect 46338 4398 46340 4450
rect 46284 4386 46340 4398
rect 46396 5124 46452 5134
rect 46396 4228 46452 5068
rect 46508 4228 46564 4238
rect 46396 4226 46564 4228
rect 46396 4174 46510 4226
rect 46562 4174 46564 4226
rect 46396 4172 46564 4174
rect 46508 4162 46564 4172
rect 46620 4114 46676 5742
rect 46732 5122 46788 6078
rect 47292 6130 47348 6188
rect 47292 6078 47294 6130
rect 47346 6078 47348 6130
rect 47292 6066 47348 6078
rect 46732 5070 46734 5122
rect 46786 5070 46788 5122
rect 46732 5058 46788 5070
rect 47180 6020 47236 6030
rect 47180 5124 47236 5964
rect 47516 5906 47572 5918
rect 47516 5854 47518 5906
rect 47570 5854 47572 5906
rect 47404 5124 47460 5134
rect 47180 5122 47460 5124
rect 47180 5070 47406 5122
rect 47458 5070 47460 5122
rect 47180 5068 47460 5070
rect 47404 5058 47460 5068
rect 47516 4340 47572 5854
rect 47740 4340 47796 4350
rect 47516 4338 47796 4340
rect 47516 4286 47742 4338
rect 47794 4286 47796 4338
rect 47516 4284 47796 4286
rect 47740 4274 47796 4284
rect 46620 4062 46622 4114
rect 46674 4062 46676 4114
rect 46620 4050 46676 4062
rect 47852 4116 47908 4126
rect 47964 4116 48020 6300
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 48076 5124 48132 5134
rect 48636 5124 48692 5134
rect 48076 5122 48692 5124
rect 48076 5070 48078 5122
rect 48130 5070 48638 5122
rect 48690 5070 48692 5122
rect 48076 5068 48692 5070
rect 48076 5058 48132 5068
rect 48636 5058 48692 5068
rect 47852 4114 48020 4116
rect 47852 4062 47854 4114
rect 47906 4062 48020 4114
rect 47852 4060 48020 4062
rect 48412 4898 48468 4910
rect 48412 4846 48414 4898
rect 48466 4846 48468 4898
rect 47852 4050 47908 4060
rect 44156 3502 44158 3554
rect 44210 3502 44212 3554
rect 44156 3490 44212 3502
rect 48412 3554 48468 4846
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 48412 3502 48414 3554
rect 48466 3502 48468 3554
rect 48412 3490 48468 3502
rect 49084 3666 49140 3678
rect 49084 3614 49086 3666
rect 49138 3614 49140 3666
rect 43708 3444 43764 3454
rect 41468 3332 41524 3342
rect 39116 3154 39172 3164
rect 41020 3330 41524 3332
rect 41020 3278 41470 3330
rect 41522 3278 41524 3330
rect 41020 3276 41524 3278
rect 39004 1474 39060 1484
rect 7868 1362 7924 1372
rect 41020 800 41076 3276
rect 41468 3266 41524 3276
rect 43708 800 43764 3388
rect 44940 3444 44996 3454
rect 49084 3388 49140 3614
rect 44940 3330 44996 3388
rect 44940 3278 44942 3330
rect 44994 3278 44996 3330
rect 44940 3266 44996 3278
rect 48524 3332 49140 3388
rect 51772 3668 51828 3678
rect 48524 1652 48580 3332
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 48412 1596 48580 1652
rect 48412 800 48468 1596
rect 51772 800 51828 3612
rect 52108 3554 52164 6412
rect 58156 5682 58212 5694
rect 58156 5630 58158 5682
rect 58210 5630 58212 5682
rect 58156 5460 58212 5630
rect 58156 5394 58212 5404
rect 58156 5234 58212 5246
rect 58156 5182 58158 5234
rect 58210 5182 58212 5234
rect 58156 4788 58212 5182
rect 58156 4722 58212 4732
rect 58156 4450 58212 4462
rect 58156 4398 58158 4450
rect 58210 4398 58212 4450
rect 58156 4116 58212 4398
rect 58156 4050 58212 4060
rect 52892 3668 52948 3678
rect 52892 3574 52948 3612
rect 52108 3502 52110 3554
rect 52162 3502 52164 3554
rect 52108 3490 52164 3502
rect 57708 3330 57764 3342
rect 57708 3278 57710 3330
rect 57762 3278 57764 3330
rect 57708 2772 57764 3278
rect 58156 3332 58212 3342
rect 58156 3238 58212 3276
rect 57708 2706 57764 2716
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 40992 0 41104 800
rect 43680 0 43792 800
rect 48384 0 48496 800
rect 51744 0 51856 800
<< via2 >>
rect 15372 57148 15428 57204
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 1708 53788 1764 53844
rect 14924 53452 14980 53508
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 14140 52220 14196 52276
rect 11900 51100 11956 51156
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 8204 46508 8260 46564
rect 11228 49532 11284 49588
rect 11676 49698 11732 49700
rect 11676 49646 11678 49698
rect 11678 49646 11730 49698
rect 11730 49646 11732 49698
rect 11676 49644 11732 49646
rect 11228 46562 11284 46564
rect 11228 46510 11230 46562
rect 11230 46510 11282 46562
rect 11282 46510 11284 46562
rect 11228 46508 11284 46510
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 8092 45164 8148 45220
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 1708 41298 1764 41300
rect 1708 41246 1710 41298
rect 1710 41246 1762 41298
rect 1762 41246 1764 41298
rect 1708 41244 1764 41246
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 1708 37826 1764 37828
rect 1708 37774 1710 37826
rect 1710 37774 1762 37826
rect 1762 37774 1764 37826
rect 1708 37772 1764 37774
rect 7868 37266 7924 37268
rect 7868 37214 7870 37266
rect 7870 37214 7922 37266
rect 7922 37214 7924 37266
rect 7868 37212 7924 37214
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 8092 34636 8148 34692
rect 4172 34130 4228 34132
rect 4172 34078 4174 34130
rect 4174 34078 4226 34130
rect 4226 34078 4228 34130
rect 4172 34076 4228 34078
rect 4844 34076 4900 34132
rect 1932 33906 1988 33908
rect 1932 33854 1934 33906
rect 1934 33854 1986 33906
rect 1986 33854 1988 33906
rect 1932 33852 1988 33854
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4844 33628 4900 33684
rect 4284 33346 4340 33348
rect 4284 33294 4286 33346
rect 4286 33294 4338 33346
rect 4338 33294 4340 33346
rect 4284 33292 4340 33294
rect 1932 32956 1988 33012
rect 1708 32284 1764 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 9884 46396 9940 46452
rect 8876 41692 8932 41748
rect 10556 45330 10612 45332
rect 10556 45278 10558 45330
rect 10558 45278 10610 45330
rect 10610 45278 10612 45330
rect 10556 45276 10612 45278
rect 10108 44322 10164 44324
rect 10108 44270 10110 44322
rect 10110 44270 10162 44322
rect 10162 44270 10164 44322
rect 10108 44268 10164 44270
rect 9996 43484 10052 43540
rect 10332 44098 10388 44100
rect 10332 44046 10334 44098
rect 10334 44046 10386 44098
rect 10386 44046 10388 44098
rect 10332 44044 10388 44046
rect 10444 43820 10500 43876
rect 10444 43538 10500 43540
rect 10444 43486 10446 43538
rect 10446 43486 10498 43538
rect 10498 43486 10500 43538
rect 10444 43484 10500 43486
rect 10220 41298 10276 41300
rect 10220 41246 10222 41298
rect 10222 41246 10274 41298
rect 10274 41246 10276 41298
rect 10220 41244 10276 41246
rect 9660 41132 9716 41188
rect 8764 40962 8820 40964
rect 8764 40910 8766 40962
rect 8766 40910 8818 40962
rect 8818 40910 8820 40962
rect 8764 40908 8820 40910
rect 8764 39564 8820 39620
rect 9772 40908 9828 40964
rect 9772 40348 9828 40404
rect 9436 39618 9492 39620
rect 9436 39566 9438 39618
rect 9438 39566 9490 39618
rect 9490 39566 9492 39618
rect 9436 39564 9492 39566
rect 8988 37548 9044 37604
rect 8316 35756 8372 35812
rect 8988 34914 9044 34916
rect 8988 34862 8990 34914
rect 8990 34862 9042 34914
rect 9042 34862 9044 34914
rect 8988 34860 9044 34862
rect 12012 50652 12068 50708
rect 12908 50706 12964 50708
rect 12908 50654 12910 50706
rect 12910 50654 12962 50706
rect 12962 50654 12964 50706
rect 12908 50652 12964 50654
rect 13468 50652 13524 50708
rect 14364 50988 14420 51044
rect 12124 49698 12180 49700
rect 12124 49646 12126 49698
rect 12126 49646 12178 49698
rect 12178 49646 12180 49698
rect 12124 49644 12180 49646
rect 12460 49644 12516 49700
rect 12012 49586 12068 49588
rect 12012 49534 12014 49586
rect 12014 49534 12066 49586
rect 12066 49534 12068 49586
rect 12012 49532 12068 49534
rect 13468 49698 13524 49700
rect 13468 49646 13470 49698
rect 13470 49646 13522 49698
rect 13522 49646 13524 49698
rect 13468 49644 13524 49646
rect 12460 47180 12516 47236
rect 12460 46396 12516 46452
rect 12348 46060 12404 46116
rect 11116 44994 11172 44996
rect 11116 44942 11118 44994
rect 11118 44942 11170 44994
rect 11170 44942 11172 44994
rect 11116 44940 11172 44942
rect 10892 44322 10948 44324
rect 10892 44270 10894 44322
rect 10894 44270 10946 44322
rect 10946 44270 10948 44322
rect 10892 44268 10948 44270
rect 10780 43484 10836 43540
rect 11228 43820 11284 43876
rect 10892 43314 10948 43316
rect 10892 43262 10894 43314
rect 10894 43262 10946 43314
rect 10946 43262 10948 43314
rect 10892 43260 10948 43262
rect 11564 43260 11620 43316
rect 12460 46002 12516 46004
rect 12460 45950 12462 46002
rect 12462 45950 12514 46002
rect 12514 45950 12516 46002
rect 12460 45948 12516 45950
rect 12012 44268 12068 44324
rect 11004 41244 11060 41300
rect 10668 40572 10724 40628
rect 10332 38780 10388 38836
rect 11004 40402 11060 40404
rect 11004 40350 11006 40402
rect 11006 40350 11058 40402
rect 11058 40350 11060 40402
rect 11004 40348 11060 40350
rect 11340 40348 11396 40404
rect 11564 39676 11620 39732
rect 9660 37884 9716 37940
rect 10444 37884 10500 37940
rect 11452 39340 11508 39396
rect 10556 37212 10612 37268
rect 9660 37100 9716 37156
rect 10108 36876 10164 36932
rect 9324 36316 9380 36372
rect 9212 36258 9268 36260
rect 9212 36206 9214 36258
rect 9214 36206 9266 36258
rect 9266 36206 9268 36258
rect 9212 36204 9268 36206
rect 9996 36370 10052 36372
rect 9996 36318 9998 36370
rect 9998 36318 10050 36370
rect 10050 36318 10052 36370
rect 9996 36316 10052 36318
rect 9548 35810 9604 35812
rect 9548 35758 9550 35810
rect 9550 35758 9602 35810
rect 9602 35758 9604 35810
rect 9548 35756 9604 35758
rect 8540 34188 8596 34244
rect 9996 34860 10052 34916
rect 1932 31890 1988 31892
rect 1932 31838 1934 31890
rect 1934 31838 1986 31890
rect 1986 31838 1988 31890
rect 1932 31836 1988 31838
rect 1932 30882 1988 30884
rect 1932 30830 1934 30882
rect 1934 30830 1986 30882
rect 1986 30830 1988 30882
rect 1932 30828 1988 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4284 30380 4340 30436
rect 1708 30322 1764 30324
rect 1708 30270 1710 30322
rect 1710 30270 1762 30322
rect 1762 30270 1764 30322
rect 1708 30268 1764 30270
rect 2156 29596 2212 29652
rect 4284 29484 4340 29540
rect 1932 29202 1988 29204
rect 1932 29150 1934 29202
rect 1934 29150 1986 29202
rect 1986 29150 1988 29202
rect 1932 29148 1988 29150
rect 4956 29148 5012 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6076 30994 6132 30996
rect 6076 30942 6078 30994
rect 6078 30942 6130 30994
rect 6130 30942 6132 30994
rect 6076 30940 6132 30942
rect 8876 33292 8932 33348
rect 8876 32508 8932 32564
rect 8988 31724 9044 31780
rect 8764 31612 8820 31668
rect 11340 39004 11396 39060
rect 10892 38946 10948 38948
rect 10892 38894 10894 38946
rect 10894 38894 10946 38946
rect 10946 38894 10948 38946
rect 10892 38892 10948 38894
rect 11116 37938 11172 37940
rect 11116 37886 11118 37938
rect 11118 37886 11170 37938
rect 11170 37886 11172 37938
rect 11116 37884 11172 37886
rect 10892 37266 10948 37268
rect 10892 37214 10894 37266
rect 10894 37214 10946 37266
rect 10946 37214 10948 37266
rect 10892 37212 10948 37214
rect 11004 36316 11060 36372
rect 10444 34188 10500 34244
rect 9996 33346 10052 33348
rect 9996 33294 9998 33346
rect 9998 33294 10050 33346
rect 10050 33294 10052 33346
rect 9996 33292 10052 33294
rect 10892 35644 10948 35700
rect 10780 35026 10836 35028
rect 10780 34974 10782 35026
rect 10782 34974 10834 35026
rect 10834 34974 10836 35026
rect 10780 34972 10836 34974
rect 10668 34242 10724 34244
rect 10668 34190 10670 34242
rect 10670 34190 10722 34242
rect 10722 34190 10724 34242
rect 10668 34188 10724 34190
rect 10892 34076 10948 34132
rect 10780 33346 10836 33348
rect 10780 33294 10782 33346
rect 10782 33294 10834 33346
rect 10834 33294 10836 33346
rect 10780 33292 10836 33294
rect 10556 33180 10612 33236
rect 11228 37100 11284 37156
rect 11452 38780 11508 38836
rect 11452 36876 11508 36932
rect 11452 36258 11508 36260
rect 11452 36206 11454 36258
rect 11454 36206 11506 36258
rect 11506 36206 11508 36258
rect 11452 36204 11508 36206
rect 11340 35810 11396 35812
rect 11340 35758 11342 35810
rect 11342 35758 11394 35810
rect 11394 35758 11396 35810
rect 11340 35756 11396 35758
rect 10220 32508 10276 32564
rect 10668 32562 10724 32564
rect 10668 32510 10670 32562
rect 10670 32510 10722 32562
rect 10722 32510 10724 32562
rect 10668 32508 10724 32510
rect 11228 32844 11284 32900
rect 13804 49196 13860 49252
rect 13580 48972 13636 49028
rect 13356 48242 13412 48244
rect 13356 48190 13358 48242
rect 13358 48190 13410 48242
rect 13410 48190 13412 48242
rect 13356 48188 13412 48190
rect 14028 49586 14084 49588
rect 14028 49534 14030 49586
rect 14030 49534 14082 49586
rect 14082 49534 14084 49586
rect 14028 49532 14084 49534
rect 13916 48636 13972 48692
rect 13580 46956 13636 47012
rect 14140 48242 14196 48244
rect 14140 48190 14142 48242
rect 14142 48190 14194 48242
rect 14194 48190 14196 48242
rect 14140 48188 14196 48190
rect 12684 46450 12740 46452
rect 12684 46398 12686 46450
rect 12686 46398 12738 46450
rect 12738 46398 12740 46450
rect 12684 46396 12740 46398
rect 13020 46450 13076 46452
rect 13020 46398 13022 46450
rect 13022 46398 13074 46450
rect 13074 46398 13076 46450
rect 13020 46396 13076 46398
rect 12572 43932 12628 43988
rect 12796 45500 12852 45556
rect 11788 41468 11844 41524
rect 11676 39116 11732 39172
rect 12460 43484 12516 43540
rect 12460 42476 12516 42532
rect 13020 44604 13076 44660
rect 13468 45612 13524 45668
rect 13692 46114 13748 46116
rect 13692 46062 13694 46114
rect 13694 46062 13746 46114
rect 13746 46062 13748 46114
rect 13692 46060 13748 46062
rect 13692 44604 13748 44660
rect 14588 50482 14644 50484
rect 14588 50430 14590 50482
rect 14590 50430 14642 50482
rect 14642 50430 14644 50482
rect 14588 50428 14644 50430
rect 14588 49420 14644 49476
rect 14700 49698 14756 49700
rect 14700 49646 14702 49698
rect 14702 49646 14754 49698
rect 14754 49646 14756 49698
rect 14700 49644 14756 49646
rect 14476 49308 14532 49364
rect 14028 45948 14084 46004
rect 14140 46396 14196 46452
rect 14812 49196 14868 49252
rect 14588 46060 14644 46116
rect 14364 45948 14420 46004
rect 14252 45890 14308 45892
rect 14252 45838 14254 45890
rect 14254 45838 14306 45890
rect 14306 45838 14308 45890
rect 14252 45836 14308 45838
rect 14252 45612 14308 45668
rect 14140 44492 14196 44548
rect 13020 43260 13076 43316
rect 13692 43314 13748 43316
rect 13692 43262 13694 43314
rect 13694 43262 13746 43314
rect 13746 43262 13748 43314
rect 13692 43260 13748 43262
rect 13580 42476 13636 42532
rect 13244 42028 13300 42084
rect 12684 41468 12740 41524
rect 12348 41186 12404 41188
rect 12348 41134 12350 41186
rect 12350 41134 12402 41186
rect 12402 41134 12404 41186
rect 12348 41132 12404 41134
rect 12684 41074 12740 41076
rect 12684 41022 12686 41074
rect 12686 41022 12738 41074
rect 12738 41022 12740 41074
rect 12684 41020 12740 41022
rect 12012 40962 12068 40964
rect 12012 40910 12014 40962
rect 12014 40910 12066 40962
rect 12066 40910 12068 40962
rect 12012 40908 12068 40910
rect 12012 40684 12068 40740
rect 12684 40236 12740 40292
rect 13468 40684 13524 40740
rect 13356 40572 13412 40628
rect 13244 40514 13300 40516
rect 13244 40462 13246 40514
rect 13246 40462 13298 40514
rect 13298 40462 13300 40514
rect 13244 40460 13300 40462
rect 13916 41970 13972 41972
rect 13916 41918 13918 41970
rect 13918 41918 13970 41970
rect 13970 41918 13972 41970
rect 13916 41916 13972 41918
rect 13468 40236 13524 40292
rect 12908 39618 12964 39620
rect 12908 39566 12910 39618
rect 12910 39566 12962 39618
rect 12962 39566 12964 39618
rect 12908 39564 12964 39566
rect 13580 39564 13636 39620
rect 12460 39394 12516 39396
rect 12460 39342 12462 39394
rect 12462 39342 12514 39394
rect 12514 39342 12516 39394
rect 12460 39340 12516 39342
rect 13804 39340 13860 39396
rect 11788 38780 11844 38836
rect 11900 38668 11956 38724
rect 13468 38834 13524 38836
rect 13468 38782 13470 38834
rect 13470 38782 13522 38834
rect 13522 38782 13524 38834
rect 13468 38780 13524 38782
rect 13244 38722 13300 38724
rect 13244 38670 13246 38722
rect 13246 38670 13298 38722
rect 13298 38670 13300 38722
rect 13244 38668 13300 38670
rect 12908 38162 12964 38164
rect 12908 38110 12910 38162
rect 12910 38110 12962 38162
rect 12962 38110 12964 38162
rect 12908 38108 12964 38110
rect 12124 37436 12180 37492
rect 11676 35810 11732 35812
rect 11676 35758 11678 35810
rect 11678 35758 11730 35810
rect 11730 35758 11732 35810
rect 11676 35756 11732 35758
rect 12460 36428 12516 36484
rect 12348 35756 12404 35812
rect 12572 36316 12628 36372
rect 11900 35698 11956 35700
rect 11900 35646 11902 35698
rect 11902 35646 11954 35698
rect 11954 35646 11956 35698
rect 11900 35644 11956 35646
rect 11564 34972 11620 35028
rect 11116 32060 11172 32116
rect 11788 35532 11844 35588
rect 12236 34748 12292 34804
rect 11676 33628 11732 33684
rect 12572 34636 12628 34692
rect 12796 37266 12852 37268
rect 12796 37214 12798 37266
rect 12798 37214 12850 37266
rect 12850 37214 12852 37266
rect 12796 37212 12852 37214
rect 12684 33346 12740 33348
rect 12684 33294 12686 33346
rect 12686 33294 12738 33346
rect 12738 33294 12740 33346
rect 12684 33292 12740 33294
rect 12124 33068 12180 33124
rect 10556 31890 10612 31892
rect 10556 31838 10558 31890
rect 10558 31838 10610 31890
rect 10610 31838 10612 31890
rect 10556 31836 10612 31838
rect 11788 32508 11844 32564
rect 9996 31778 10052 31780
rect 9996 31726 9998 31778
rect 9998 31726 10050 31778
rect 10050 31726 10052 31778
rect 9996 31724 10052 31726
rect 10892 31778 10948 31780
rect 10892 31726 10894 31778
rect 10894 31726 10946 31778
rect 10946 31726 10948 31778
rect 10892 31724 10948 31726
rect 12460 32562 12516 32564
rect 12460 32510 12462 32562
rect 12462 32510 12514 32562
rect 12514 32510 12516 32562
rect 12460 32508 12516 32510
rect 12908 37042 12964 37044
rect 12908 36990 12910 37042
rect 12910 36990 12962 37042
rect 12962 36990 12964 37042
rect 12908 36988 12964 36990
rect 13244 36316 13300 36372
rect 12908 35196 12964 35252
rect 12908 34748 12964 34804
rect 13804 38050 13860 38052
rect 13804 37998 13806 38050
rect 13806 37998 13858 38050
rect 13858 37998 13860 38050
rect 13804 37996 13860 37998
rect 14028 39004 14084 39060
rect 13916 38108 13972 38164
rect 14028 38050 14084 38052
rect 14028 37998 14030 38050
rect 14030 37998 14082 38050
rect 14082 37998 14084 38050
rect 14028 37996 14084 37998
rect 14364 45276 14420 45332
rect 14476 44994 14532 44996
rect 14476 44942 14478 44994
rect 14478 44942 14530 44994
rect 14530 44942 14532 44994
rect 14476 44940 14532 44942
rect 15260 50482 15316 50484
rect 15260 50430 15262 50482
rect 15262 50430 15314 50482
rect 15314 50430 15316 50482
rect 15260 50428 15316 50430
rect 15148 50316 15204 50372
rect 15260 49756 15316 49812
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 18060 55692 18116 55748
rect 17836 54684 17892 54740
rect 16044 53618 16100 53620
rect 16044 53566 16046 53618
rect 16046 53566 16098 53618
rect 16098 53566 16100 53618
rect 16044 53564 16100 53566
rect 15596 52722 15652 52724
rect 15596 52670 15598 52722
rect 15598 52670 15650 52722
rect 15650 52670 15652 52722
rect 15596 52668 15652 52670
rect 15484 51548 15540 51604
rect 15484 51212 15540 51268
rect 15708 50876 15764 50932
rect 16492 53506 16548 53508
rect 16492 53454 16494 53506
rect 16494 53454 16546 53506
rect 16546 53454 16548 53506
rect 16492 53452 16548 53454
rect 16940 53788 16996 53844
rect 17836 53788 17892 53844
rect 16716 53618 16772 53620
rect 16716 53566 16718 53618
rect 16718 53566 16770 53618
rect 16770 53566 16772 53618
rect 16716 53564 16772 53566
rect 17500 53506 17556 53508
rect 17500 53454 17502 53506
rect 17502 53454 17554 53506
rect 17554 53454 17556 53506
rect 17500 53452 17556 53454
rect 17164 53228 17220 53284
rect 17724 53116 17780 53172
rect 17500 53058 17556 53060
rect 17500 53006 17502 53058
rect 17502 53006 17554 53058
rect 17554 53006 17556 53058
rect 17500 53004 17556 53006
rect 17612 52946 17668 52948
rect 17612 52894 17614 52946
rect 17614 52894 17666 52946
rect 17666 52894 17668 52946
rect 17612 52892 17668 52894
rect 16940 52556 16996 52612
rect 17164 51996 17220 52052
rect 16716 51548 16772 51604
rect 16268 51378 16324 51380
rect 16268 51326 16270 51378
rect 16270 51326 16322 51378
rect 16322 51326 16324 51378
rect 16268 51324 16324 51326
rect 15596 50540 15652 50596
rect 15484 50204 15540 50260
rect 15036 46786 15092 46788
rect 15036 46734 15038 46786
rect 15038 46734 15090 46786
rect 15090 46734 15092 46786
rect 15036 46732 15092 46734
rect 14924 45890 14980 45892
rect 14924 45838 14926 45890
rect 14926 45838 14978 45890
rect 14978 45838 14980 45890
rect 14924 45836 14980 45838
rect 14812 45612 14868 45668
rect 14924 45276 14980 45332
rect 14364 44434 14420 44436
rect 14364 44382 14366 44434
rect 14366 44382 14418 44434
rect 14418 44382 14420 44434
rect 14364 44380 14420 44382
rect 14252 40124 14308 40180
rect 15036 44492 15092 44548
rect 14588 44380 14644 44436
rect 14588 42028 14644 42084
rect 14476 41692 14532 41748
rect 14812 41356 14868 41412
rect 15372 48076 15428 48132
rect 15708 50370 15764 50372
rect 15708 50318 15710 50370
rect 15710 50318 15762 50370
rect 15762 50318 15764 50370
rect 15708 50316 15764 50318
rect 15708 48076 15764 48132
rect 15596 47234 15652 47236
rect 15596 47182 15598 47234
rect 15598 47182 15650 47234
rect 15650 47182 15652 47234
rect 15596 47180 15652 47182
rect 15596 45836 15652 45892
rect 15484 45388 15540 45444
rect 15596 45612 15652 45668
rect 15372 45164 15428 45220
rect 15372 44380 15428 44436
rect 16380 51266 16436 51268
rect 16380 51214 16382 51266
rect 16382 51214 16434 51266
rect 16434 51214 16436 51266
rect 16380 51212 16436 51214
rect 17500 51266 17556 51268
rect 17500 51214 17502 51266
rect 17502 51214 17554 51266
rect 17554 51214 17556 51266
rect 17500 51212 17556 51214
rect 18732 55074 18788 55076
rect 18732 55022 18734 55074
rect 18734 55022 18786 55074
rect 18786 55022 18788 55074
rect 18732 55020 18788 55022
rect 19180 55074 19236 55076
rect 19180 55022 19182 55074
rect 19182 55022 19234 55074
rect 19234 55022 19236 55074
rect 19180 55020 19236 55022
rect 19068 54402 19124 54404
rect 19068 54350 19070 54402
rect 19070 54350 19122 54402
rect 19122 54350 19124 54402
rect 19068 54348 19124 54350
rect 18844 53228 18900 53284
rect 18620 53058 18676 53060
rect 18620 53006 18622 53058
rect 18622 53006 18674 53058
rect 18674 53006 18676 53058
rect 18620 53004 18676 53006
rect 18172 52556 18228 52612
rect 18396 52780 18452 52836
rect 18060 52108 18116 52164
rect 17388 50706 17444 50708
rect 17388 50654 17390 50706
rect 17390 50654 17442 50706
rect 17442 50654 17444 50706
rect 17388 50652 17444 50654
rect 18284 52220 18340 52276
rect 16716 50092 16772 50148
rect 16156 48636 16212 48692
rect 16380 49756 16436 49812
rect 16828 49698 16884 49700
rect 16828 49646 16830 49698
rect 16830 49646 16882 49698
rect 16882 49646 16884 49698
rect 16828 49644 16884 49646
rect 17052 50092 17108 50148
rect 17836 49922 17892 49924
rect 17836 49870 17838 49922
rect 17838 49870 17890 49922
rect 17890 49870 17892 49922
rect 17836 49868 17892 49870
rect 18284 51212 18340 51268
rect 17500 49810 17556 49812
rect 17500 49758 17502 49810
rect 17502 49758 17554 49810
rect 17554 49758 17556 49810
rect 17500 49756 17556 49758
rect 16940 49308 16996 49364
rect 17836 49308 17892 49364
rect 16604 49026 16660 49028
rect 16604 48974 16606 49026
rect 16606 48974 16658 49026
rect 16658 48974 16660 49026
rect 16604 48972 16660 48974
rect 16268 48130 16324 48132
rect 16268 48078 16270 48130
rect 16270 48078 16322 48130
rect 16322 48078 16324 48130
rect 16268 48076 16324 48078
rect 16604 48748 16660 48804
rect 16716 47404 16772 47460
rect 16044 46956 16100 47012
rect 16604 46956 16660 47012
rect 16268 46562 16324 46564
rect 16268 46510 16270 46562
rect 16270 46510 16322 46562
rect 16322 46510 16324 46562
rect 16268 46508 16324 46510
rect 16492 46450 16548 46452
rect 16492 46398 16494 46450
rect 16494 46398 16546 46450
rect 16546 46398 16548 46450
rect 16492 46396 16548 46398
rect 15820 44546 15876 44548
rect 15820 44494 15822 44546
rect 15822 44494 15874 44546
rect 15874 44494 15876 44546
rect 15820 44492 15876 44494
rect 16044 45724 16100 45780
rect 15708 43538 15764 43540
rect 15708 43486 15710 43538
rect 15710 43486 15762 43538
rect 15762 43486 15764 43538
rect 15708 43484 15764 43486
rect 15932 44322 15988 44324
rect 15932 44270 15934 44322
rect 15934 44270 15986 44322
rect 15986 44270 15988 44322
rect 15932 44268 15988 44270
rect 16268 45890 16324 45892
rect 16268 45838 16270 45890
rect 16270 45838 16322 45890
rect 16322 45838 16324 45890
rect 16268 45836 16324 45838
rect 16828 46898 16884 46900
rect 16828 46846 16830 46898
rect 16830 46846 16882 46898
rect 16882 46846 16884 46898
rect 16828 46844 16884 46846
rect 16716 46172 16772 46228
rect 16828 45948 16884 46004
rect 16940 45890 16996 45892
rect 16940 45838 16942 45890
rect 16942 45838 16994 45890
rect 16994 45838 16996 45890
rect 16940 45836 16996 45838
rect 16492 45500 16548 45556
rect 16716 45218 16772 45220
rect 16716 45166 16718 45218
rect 16718 45166 16770 45218
rect 16770 45166 16772 45218
rect 16716 45164 16772 45166
rect 16268 44940 16324 44996
rect 16940 44828 16996 44884
rect 16268 44380 16324 44436
rect 16716 44380 16772 44436
rect 16492 44098 16548 44100
rect 16492 44046 16494 44098
rect 16494 44046 16546 44098
rect 16546 44046 16548 44098
rect 16492 44044 16548 44046
rect 16268 43708 16324 43764
rect 16156 43596 16212 43652
rect 16380 43650 16436 43652
rect 16380 43598 16382 43650
rect 16382 43598 16434 43650
rect 16434 43598 16436 43650
rect 16380 43596 16436 43598
rect 16604 43596 16660 43652
rect 15484 43260 15540 43316
rect 15260 42140 15316 42196
rect 15036 42028 15092 42084
rect 15260 41916 15316 41972
rect 15260 41746 15316 41748
rect 15260 41694 15262 41746
rect 15262 41694 15314 41746
rect 15314 41694 15316 41746
rect 15260 41692 15316 41694
rect 15148 41580 15204 41636
rect 14588 41244 14644 41300
rect 14476 40012 14532 40068
rect 14476 39730 14532 39732
rect 14476 39678 14478 39730
rect 14478 39678 14530 39730
rect 14530 39678 14532 39730
rect 14476 39676 14532 39678
rect 14364 39340 14420 39396
rect 14812 40236 14868 40292
rect 15260 41298 15316 41300
rect 15260 41246 15262 41298
rect 15262 41246 15314 41298
rect 15314 41246 15316 41298
rect 15260 41244 15316 41246
rect 15148 40460 15204 40516
rect 15036 40348 15092 40404
rect 14812 39004 14868 39060
rect 15148 38946 15204 38948
rect 15148 38894 15150 38946
rect 15150 38894 15202 38946
rect 15202 38894 15204 38946
rect 15148 38892 15204 38894
rect 14700 38332 14756 38388
rect 14252 37324 14308 37380
rect 14140 36428 14196 36484
rect 13692 35756 13748 35812
rect 14028 35532 14084 35588
rect 13356 33068 13412 33124
rect 13468 35196 13524 35252
rect 13580 34690 13636 34692
rect 13580 34638 13582 34690
rect 13582 34638 13634 34690
rect 13634 34638 13636 34690
rect 13580 34636 13636 34638
rect 13580 34130 13636 34132
rect 13580 34078 13582 34130
rect 13582 34078 13634 34130
rect 13634 34078 13636 34130
rect 13580 34076 13636 34078
rect 13692 33740 13748 33796
rect 14252 33180 14308 33236
rect 13468 32396 13524 32452
rect 13580 32674 13636 32676
rect 13580 32622 13582 32674
rect 13582 32622 13634 32674
rect 13634 32622 13636 32674
rect 13580 32620 13636 32622
rect 12796 31948 12852 32004
rect 14028 32562 14084 32564
rect 14028 32510 14030 32562
rect 14030 32510 14082 32562
rect 14082 32510 14084 32562
rect 14028 32508 14084 32510
rect 14140 32396 14196 32452
rect 9884 31164 9940 31220
rect 12348 31218 12404 31220
rect 12348 31166 12350 31218
rect 12350 31166 12402 31218
rect 12402 31166 12404 31218
rect 12348 31164 12404 31166
rect 14588 35922 14644 35924
rect 14588 35870 14590 35922
rect 14590 35870 14642 35922
rect 14642 35870 14644 35922
rect 14588 35868 14644 35870
rect 14588 35532 14644 35588
rect 14700 35196 14756 35252
rect 14476 33404 14532 33460
rect 14588 33852 14644 33908
rect 14924 34860 14980 34916
rect 15036 34748 15092 34804
rect 15596 42588 15652 42644
rect 16380 43260 16436 43316
rect 16156 42140 16212 42196
rect 15708 41916 15764 41972
rect 16044 41970 16100 41972
rect 16044 41918 16046 41970
rect 16046 41918 16098 41970
rect 16098 41918 16100 41970
rect 16044 41916 16100 41918
rect 16156 41468 16212 41524
rect 15708 40684 15764 40740
rect 15484 40348 15540 40404
rect 15596 40290 15652 40292
rect 15596 40238 15598 40290
rect 15598 40238 15650 40290
rect 15650 40238 15652 40290
rect 15596 40236 15652 40238
rect 16268 40514 16324 40516
rect 16268 40462 16270 40514
rect 16270 40462 16322 40514
rect 16322 40462 16324 40514
rect 16268 40460 16324 40462
rect 17052 44492 17108 44548
rect 17164 48076 17220 48132
rect 17052 44268 17108 44324
rect 18396 51100 18452 51156
rect 18396 50764 18452 50820
rect 19964 55186 20020 55188
rect 19964 55134 19966 55186
rect 19966 55134 20018 55186
rect 20018 55134 20020 55186
rect 19964 55132 20020 55134
rect 19852 55074 19908 55076
rect 19852 55022 19854 55074
rect 19854 55022 19906 55074
rect 19906 55022 19908 55074
rect 19852 55020 19908 55022
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 20412 54514 20468 54516
rect 20412 54462 20414 54514
rect 20414 54462 20466 54514
rect 20466 54462 20468 54514
rect 20412 54460 20468 54462
rect 19852 54236 19908 54292
rect 19740 53842 19796 53844
rect 19740 53790 19742 53842
rect 19742 53790 19794 53842
rect 19794 53790 19796 53842
rect 19740 53788 19796 53790
rect 19628 53676 19684 53732
rect 20860 54012 20916 54068
rect 21196 54348 21252 54404
rect 20300 53676 20356 53732
rect 19292 53116 19348 53172
rect 18844 51324 18900 51380
rect 19068 52892 19124 52948
rect 19628 53228 19684 53284
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19852 52780 19908 52836
rect 19180 52556 19236 52612
rect 19964 52556 20020 52612
rect 19180 52108 19236 52164
rect 19404 52220 19460 52276
rect 19628 51772 19684 51828
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19180 51324 19236 51380
rect 19292 51212 19348 51268
rect 18732 50988 18788 51044
rect 18956 50092 19012 50148
rect 18620 49868 18676 49924
rect 18956 49644 19012 49700
rect 18396 49084 18452 49140
rect 19068 49084 19124 49140
rect 18956 49026 19012 49028
rect 18956 48974 18958 49026
rect 18958 48974 19010 49026
rect 19010 48974 19012 49026
rect 18956 48972 19012 48974
rect 18508 48130 18564 48132
rect 18508 48078 18510 48130
rect 18510 48078 18562 48130
rect 18562 48078 18564 48130
rect 18508 48076 18564 48078
rect 17948 47740 18004 47796
rect 17836 47292 17892 47348
rect 17500 47180 17556 47236
rect 17388 46450 17444 46452
rect 17388 46398 17390 46450
rect 17390 46398 17442 46450
rect 17442 46398 17444 46450
rect 17388 46396 17444 46398
rect 17500 45948 17556 46004
rect 19628 50988 19684 51044
rect 19516 50652 19572 50708
rect 19628 50764 19684 50820
rect 20188 51100 20244 51156
rect 19404 49980 19460 50036
rect 20412 53506 20468 53508
rect 20412 53454 20414 53506
rect 20414 53454 20466 53506
rect 20466 53454 20468 53506
rect 20412 53452 20468 53454
rect 20524 53228 20580 53284
rect 20748 53506 20804 53508
rect 20748 53454 20750 53506
rect 20750 53454 20802 53506
rect 20802 53454 20804 53506
rect 20748 53452 20804 53454
rect 20524 52444 20580 52500
rect 20636 52332 20692 52388
rect 20524 52050 20580 52052
rect 20524 51998 20526 52050
rect 20526 51998 20578 52050
rect 20578 51998 20580 52050
rect 20524 51996 20580 51998
rect 20860 52162 20916 52164
rect 20860 52110 20862 52162
rect 20862 52110 20914 52162
rect 20914 52110 20916 52162
rect 20860 52108 20916 52110
rect 22204 54796 22260 54852
rect 21644 54572 21700 54628
rect 21308 54236 21364 54292
rect 21420 54460 21476 54516
rect 22764 54796 22820 54852
rect 22204 54514 22260 54516
rect 22204 54462 22206 54514
rect 22206 54462 22258 54514
rect 22258 54462 22260 54514
rect 22204 54460 22260 54462
rect 22428 54572 22484 54628
rect 21532 54348 21588 54404
rect 21196 52834 21252 52836
rect 21196 52782 21198 52834
rect 21198 52782 21250 52834
rect 21250 52782 21252 52834
rect 21196 52780 21252 52782
rect 21420 52332 21476 52388
rect 20300 50316 20356 50372
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19628 49922 19684 49924
rect 19628 49870 19630 49922
rect 19630 49870 19682 49922
rect 19682 49870 19684 49922
rect 19628 49868 19684 49870
rect 19292 49196 19348 49252
rect 19292 48860 19348 48916
rect 18844 47740 18900 47796
rect 17948 46956 18004 47012
rect 18060 46786 18116 46788
rect 18060 46734 18062 46786
rect 18062 46734 18114 46786
rect 18114 46734 18116 46786
rect 18060 46732 18116 46734
rect 17836 46674 17892 46676
rect 17836 46622 17838 46674
rect 17838 46622 17890 46674
rect 17890 46622 17892 46674
rect 17836 46620 17892 46622
rect 17724 46508 17780 46564
rect 17724 45890 17780 45892
rect 17724 45838 17726 45890
rect 17726 45838 17778 45890
rect 17778 45838 17780 45890
rect 17724 45836 17780 45838
rect 17388 45388 17444 45444
rect 17388 44492 17444 44548
rect 16940 43484 16996 43540
rect 16828 42812 16884 42868
rect 16604 42588 16660 42644
rect 16716 40684 16772 40740
rect 16492 40514 16548 40516
rect 16492 40462 16494 40514
rect 16494 40462 16546 40514
rect 16546 40462 16548 40514
rect 16492 40460 16548 40462
rect 16156 39004 16212 39060
rect 16044 38780 16100 38836
rect 15932 38274 15988 38276
rect 15932 38222 15934 38274
rect 15934 38222 15986 38274
rect 15986 38222 15988 38274
rect 15932 38220 15988 38222
rect 15708 38108 15764 38164
rect 16044 37996 16100 38052
rect 15820 37436 15876 37492
rect 15820 37212 15876 37268
rect 16044 37266 16100 37268
rect 16044 37214 16046 37266
rect 16046 37214 16098 37266
rect 16098 37214 16100 37266
rect 16044 37212 16100 37214
rect 15820 36482 15876 36484
rect 15820 36430 15822 36482
rect 15822 36430 15874 36482
rect 15874 36430 15876 36482
rect 15820 36428 15876 36430
rect 16044 34914 16100 34916
rect 16044 34862 16046 34914
rect 16046 34862 16098 34914
rect 16098 34862 16100 34914
rect 16044 34860 16100 34862
rect 14700 33180 14756 33236
rect 15372 33906 15428 33908
rect 15372 33854 15374 33906
rect 15374 33854 15426 33906
rect 15426 33854 15428 33906
rect 15372 33852 15428 33854
rect 15708 34354 15764 34356
rect 15708 34302 15710 34354
rect 15710 34302 15762 34354
rect 15762 34302 15764 34354
rect 15708 34300 15764 34302
rect 15596 33234 15652 33236
rect 15596 33182 15598 33234
rect 15598 33182 15650 33234
rect 15650 33182 15652 33234
rect 15596 33180 15652 33182
rect 15372 32844 15428 32900
rect 15932 32786 15988 32788
rect 15932 32734 15934 32786
rect 15934 32734 15986 32786
rect 15986 32734 15988 32786
rect 15932 32732 15988 32734
rect 14588 32508 14644 32564
rect 15148 32620 15204 32676
rect 15708 32674 15764 32676
rect 15708 32622 15710 32674
rect 15710 32622 15762 32674
rect 15762 32622 15764 32674
rect 15708 32620 15764 32622
rect 15148 32450 15204 32452
rect 15148 32398 15150 32450
rect 15150 32398 15202 32450
rect 15202 32398 15204 32450
rect 15148 32396 15204 32398
rect 14700 31890 14756 31892
rect 14700 31838 14702 31890
rect 14702 31838 14754 31890
rect 14754 31838 14756 31890
rect 14700 31836 14756 31838
rect 14364 31500 14420 31556
rect 14700 31612 14756 31668
rect 8540 31052 8596 31108
rect 9548 31106 9604 31108
rect 9548 31054 9550 31106
rect 9550 31054 9602 31106
rect 9602 31054 9604 31106
rect 9548 31052 9604 31054
rect 9100 30380 9156 30436
rect 8316 29596 8372 29652
rect 1708 28418 1764 28420
rect 1708 28366 1710 28418
rect 1710 28366 1762 28418
rect 1762 28366 1764 28418
rect 1708 28364 1764 28366
rect 2044 28082 2100 28084
rect 2044 28030 2046 28082
rect 2046 28030 2098 28082
rect 2098 28030 2100 28082
rect 2044 28028 2100 28030
rect 6076 27858 6132 27860
rect 6076 27806 6078 27858
rect 6078 27806 6130 27858
rect 6130 27806 6132 27858
rect 6076 27804 6132 27806
rect 1708 27580 1764 27636
rect 2492 27580 2548 27636
rect 2044 27468 2100 27524
rect 1708 26908 1764 26964
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2492 26908 2548 26964
rect 1932 26236 1988 26292
rect 2268 26236 2324 26292
rect 2380 26124 2436 26180
rect 2380 25564 2436 25620
rect 2716 26514 2772 26516
rect 2716 26462 2718 26514
rect 2718 26462 2770 26514
rect 2770 26462 2772 26514
rect 2716 26460 2772 26462
rect 3164 26178 3220 26180
rect 3164 26126 3166 26178
rect 3166 26126 3218 26178
rect 3218 26126 3220 26178
rect 3164 26124 3220 26126
rect 6300 26796 6356 26852
rect 5068 26572 5124 26628
rect 4396 26290 4452 26292
rect 4396 26238 4398 26290
rect 4398 26238 4450 26290
rect 4450 26238 4452 26290
rect 4396 26236 4452 26238
rect 4844 26290 4900 26292
rect 4844 26238 4846 26290
rect 4846 26238 4898 26290
rect 4898 26238 4900 26290
rect 4844 26236 4900 26238
rect 4284 26012 4340 26068
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1708 24892 1764 24948
rect 5740 26572 5796 26628
rect 5516 25676 5572 25732
rect 4396 25394 4452 25396
rect 4396 25342 4398 25394
rect 4398 25342 4450 25394
rect 4450 25342 4452 25394
rect 4396 25340 4452 25342
rect 5180 25340 5236 25396
rect 4172 25228 4228 25284
rect 4732 25282 4788 25284
rect 4732 25230 4734 25282
rect 4734 25230 4786 25282
rect 4786 25230 4788 25282
rect 4732 25228 4788 25230
rect 2940 24892 2996 24948
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 8876 27132 8932 27188
rect 8204 26124 8260 26180
rect 6524 25564 6580 25620
rect 6300 25228 6356 25284
rect 5964 25116 6020 25172
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 9212 27356 9268 27412
rect 8764 25676 8820 25732
rect 7980 24444 8036 24500
rect 1932 23548 1988 23604
rect 7308 23660 7364 23716
rect 4172 23324 4228 23380
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 22482 1988 22484
rect 1932 22430 1934 22482
rect 1934 22430 1986 22482
rect 1986 22430 1988 22482
rect 1932 22428 1988 22430
rect 4284 23212 4340 23268
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 6300 22204 6356 22260
rect 4284 21756 4340 21812
rect 6860 22092 6916 22148
rect 5964 21586 6020 21588
rect 5964 21534 5966 21586
rect 5966 21534 6018 21586
rect 6018 21534 6020 21586
rect 5964 21532 6020 21534
rect 1932 21474 1988 21476
rect 1932 21422 1934 21474
rect 1934 21422 1986 21474
rect 1986 21422 1988 21474
rect 1932 21420 1988 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5852 20802 5908 20804
rect 5852 20750 5854 20802
rect 5854 20750 5906 20802
rect 5906 20750 5908 20802
rect 5852 20748 5908 20750
rect 3276 20412 3332 20468
rect 1708 19010 1764 19012
rect 1708 18958 1710 19010
rect 1710 18958 1762 19010
rect 1762 18958 1764 19010
rect 1708 18956 1764 18958
rect 1708 16828 1764 16884
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 6300 20300 6356 20356
rect 6076 19906 6132 19908
rect 6076 19854 6078 19906
rect 6078 19854 6130 19906
rect 6130 19854 6132 19906
rect 6076 19852 6132 19854
rect 5740 18508 5796 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5404 17106 5460 17108
rect 5404 17054 5406 17106
rect 5406 17054 5458 17106
rect 5458 17054 5460 17106
rect 5404 17052 5460 17054
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 6076 16828 6132 16884
rect 5852 16492 5908 16548
rect 5740 15932 5796 15988
rect 5628 15314 5684 15316
rect 5628 15262 5630 15314
rect 5630 15262 5682 15314
rect 5682 15262 5684 15314
rect 5628 15260 5684 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5964 13468 6020 13524
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 6412 20018 6468 20020
rect 6412 19966 6414 20018
rect 6414 19966 6466 20018
rect 6466 19966 6468 20018
rect 6412 19964 6468 19966
rect 6748 21756 6804 21812
rect 6972 21532 7028 21588
rect 6748 19852 6804 19908
rect 6748 18562 6804 18564
rect 6748 18510 6750 18562
rect 6750 18510 6802 18562
rect 6802 18510 6804 18562
rect 6748 18508 6804 18510
rect 6524 18396 6580 18452
rect 6412 16940 6468 16996
rect 6524 15932 6580 15988
rect 6300 14700 6356 14756
rect 6188 14530 6244 14532
rect 6188 14478 6190 14530
rect 6190 14478 6242 14530
rect 6242 14478 6244 14530
rect 6188 14476 6244 14478
rect 7084 20018 7140 20020
rect 7084 19966 7086 20018
rect 7086 19966 7138 20018
rect 7138 19966 7140 20018
rect 7084 19964 7140 19966
rect 7868 23212 7924 23268
rect 7420 21756 7476 21812
rect 8764 24498 8820 24500
rect 8764 24446 8766 24498
rect 8766 24446 8818 24498
rect 8818 24446 8820 24498
rect 8764 24444 8820 24446
rect 8764 23324 8820 23380
rect 9660 27356 9716 27412
rect 12572 30380 12628 30436
rect 14588 30380 14644 30436
rect 12236 30210 12292 30212
rect 12236 30158 12238 30210
rect 12238 30158 12290 30210
rect 12290 30158 12292 30210
rect 12236 30156 12292 30158
rect 11788 29650 11844 29652
rect 11788 29598 11790 29650
rect 11790 29598 11842 29650
rect 11842 29598 11844 29650
rect 11788 29596 11844 29598
rect 12348 29596 12404 29652
rect 10108 29372 10164 29428
rect 12572 29314 12628 29316
rect 12572 29262 12574 29314
rect 12574 29262 12626 29314
rect 12626 29262 12628 29314
rect 12572 29260 12628 29262
rect 12908 28588 12964 28644
rect 10332 27186 10388 27188
rect 10332 27134 10334 27186
rect 10334 27134 10386 27186
rect 10386 27134 10388 27186
rect 10332 27132 10388 27134
rect 9436 26684 9492 26740
rect 10444 26460 10500 26516
rect 9996 26402 10052 26404
rect 9996 26350 9998 26402
rect 9998 26350 10050 26402
rect 10050 26350 10052 26402
rect 9996 26348 10052 26350
rect 11340 26684 11396 26740
rect 10780 26178 10836 26180
rect 10780 26126 10782 26178
rect 10782 26126 10834 26178
rect 10834 26126 10836 26178
rect 10780 26124 10836 26126
rect 11340 26124 11396 26180
rect 12460 26962 12516 26964
rect 12460 26910 12462 26962
rect 12462 26910 12514 26962
rect 12514 26910 12516 26962
rect 12460 26908 12516 26910
rect 13916 28642 13972 28644
rect 13916 28590 13918 28642
rect 13918 28590 13970 28642
rect 13970 28590 13972 28642
rect 13916 28588 13972 28590
rect 15596 31612 15652 31668
rect 16828 40124 16884 40180
rect 16828 39842 16884 39844
rect 16828 39790 16830 39842
rect 16830 39790 16882 39842
rect 16882 39790 16884 39842
rect 16828 39788 16884 39790
rect 16604 38892 16660 38948
rect 16828 39228 16884 39284
rect 16492 38050 16548 38052
rect 16492 37998 16494 38050
rect 16494 37998 16546 38050
rect 16546 37998 16548 38050
rect 16492 37996 16548 37998
rect 16716 36482 16772 36484
rect 16716 36430 16718 36482
rect 16718 36430 16770 36482
rect 16770 36430 16772 36482
rect 16716 36428 16772 36430
rect 17500 44156 17556 44212
rect 17948 46060 18004 46116
rect 17948 45890 18004 45892
rect 17948 45838 17950 45890
rect 17950 45838 18002 45890
rect 18002 45838 18004 45890
rect 17948 45836 18004 45838
rect 17612 44604 17668 44660
rect 17724 45052 17780 45108
rect 17836 44268 17892 44324
rect 17724 44044 17780 44100
rect 18396 47180 18452 47236
rect 18620 47180 18676 47236
rect 18508 47068 18564 47124
rect 18508 46956 18564 47012
rect 18508 46620 18564 46676
rect 18284 46172 18340 46228
rect 18508 46060 18564 46116
rect 18284 46002 18340 46004
rect 18284 45950 18286 46002
rect 18286 45950 18338 46002
rect 18338 45950 18340 46002
rect 18284 45948 18340 45950
rect 19068 47068 19124 47124
rect 18620 45836 18676 45892
rect 18732 46172 18788 46228
rect 18284 45276 18340 45332
rect 17948 44044 18004 44100
rect 17612 43650 17668 43652
rect 17612 43598 17614 43650
rect 17614 43598 17666 43650
rect 17666 43598 17668 43650
rect 17612 43596 17668 43598
rect 17724 43538 17780 43540
rect 17724 43486 17726 43538
rect 17726 43486 17778 43538
rect 17778 43486 17780 43538
rect 17724 43484 17780 43486
rect 16604 35420 16660 35476
rect 16492 34802 16548 34804
rect 16492 34750 16494 34802
rect 16494 34750 16546 34802
rect 16546 34750 16548 34802
rect 16492 34748 16548 34750
rect 16828 34636 16884 34692
rect 16492 34188 16548 34244
rect 17388 42812 17444 42868
rect 17388 42588 17444 42644
rect 17388 41916 17444 41972
rect 17164 39788 17220 39844
rect 17276 41356 17332 41412
rect 17276 41132 17332 41188
rect 17500 40348 17556 40404
rect 18172 44940 18228 44996
rect 18844 46060 18900 46116
rect 18844 45836 18900 45892
rect 18844 45612 18900 45668
rect 19292 47404 19348 47460
rect 20188 49532 20244 49588
rect 20300 48972 20356 49028
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 21308 52220 21364 52276
rect 20972 50764 21028 50820
rect 20860 50482 20916 50484
rect 20860 50430 20862 50482
rect 20862 50430 20914 50482
rect 20914 50430 20916 50482
rect 20860 50428 20916 50430
rect 20524 49532 20580 49588
rect 20748 49138 20804 49140
rect 20748 49086 20750 49138
rect 20750 49086 20802 49138
rect 20802 49086 20804 49138
rect 20748 49084 20804 49086
rect 20188 47964 20244 48020
rect 19628 47570 19684 47572
rect 19628 47518 19630 47570
rect 19630 47518 19682 47570
rect 19682 47518 19684 47570
rect 19628 47516 19684 47518
rect 19740 47346 19796 47348
rect 19740 47294 19742 47346
rect 19742 47294 19794 47346
rect 19794 47294 19796 47346
rect 19740 47292 19796 47294
rect 19404 47180 19460 47236
rect 19516 46956 19572 47012
rect 19628 47068 19684 47124
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19628 46844 19684 46900
rect 19964 46172 20020 46228
rect 20076 45890 20132 45892
rect 20076 45838 20078 45890
rect 20078 45838 20130 45890
rect 20130 45838 20132 45890
rect 20076 45836 20132 45838
rect 20300 47234 20356 47236
rect 20300 47182 20302 47234
rect 20302 47182 20354 47234
rect 20354 47182 20356 47234
rect 20300 47180 20356 47182
rect 20300 46844 20356 46900
rect 20748 48076 20804 48132
rect 20636 47404 20692 47460
rect 20524 47346 20580 47348
rect 20524 47294 20526 47346
rect 20526 47294 20578 47346
rect 20578 47294 20580 47346
rect 20524 47292 20580 47294
rect 20636 47180 20692 47236
rect 20412 46396 20468 46452
rect 21084 50034 21140 50036
rect 21084 49982 21086 50034
rect 21086 49982 21138 50034
rect 21138 49982 21140 50034
rect 21084 49980 21140 49982
rect 21420 50370 21476 50372
rect 21420 50318 21422 50370
rect 21422 50318 21474 50370
rect 21474 50318 21476 50370
rect 21420 50316 21476 50318
rect 21756 52892 21812 52948
rect 21980 52892 22036 52948
rect 21868 52162 21924 52164
rect 21868 52110 21870 52162
rect 21870 52110 21922 52162
rect 21922 52110 21924 52162
rect 21868 52108 21924 52110
rect 21756 51212 21812 51268
rect 21868 50428 21924 50484
rect 21756 49756 21812 49812
rect 21868 49084 21924 49140
rect 21644 49026 21700 49028
rect 21644 48974 21646 49026
rect 21646 48974 21698 49026
rect 21698 48974 21700 49026
rect 21644 48972 21700 48974
rect 21308 48748 21364 48804
rect 21532 48860 21588 48916
rect 21644 48466 21700 48468
rect 21644 48414 21646 48466
rect 21646 48414 21698 48466
rect 21698 48414 21700 48466
rect 21644 48412 21700 48414
rect 21196 47516 21252 47572
rect 21532 47458 21588 47460
rect 21532 47406 21534 47458
rect 21534 47406 21586 47458
rect 21586 47406 21588 47458
rect 21532 47404 21588 47406
rect 21196 47180 21252 47236
rect 20860 46172 20916 46228
rect 20636 46060 20692 46116
rect 18844 45330 18900 45332
rect 18844 45278 18846 45330
rect 18846 45278 18898 45330
rect 18898 45278 18900 45330
rect 18844 45276 18900 45278
rect 19068 45164 19124 45220
rect 18732 43708 18788 43764
rect 18732 43538 18788 43540
rect 18732 43486 18734 43538
rect 18734 43486 18786 43538
rect 18786 43486 18788 43538
rect 18732 43484 18788 43486
rect 18396 43260 18452 43316
rect 18732 43260 18788 43316
rect 19068 44268 19124 44324
rect 18172 42812 18228 42868
rect 18284 42700 18340 42756
rect 18844 42700 18900 42756
rect 18284 42252 18340 42308
rect 18732 42252 18788 42308
rect 18956 42252 19012 42308
rect 19068 42700 19124 42756
rect 19516 45666 19572 45668
rect 19516 45614 19518 45666
rect 19518 45614 19570 45666
rect 19570 45614 19572 45666
rect 19516 45612 19572 45614
rect 20300 45666 20356 45668
rect 20300 45614 20302 45666
rect 20302 45614 20354 45666
rect 20354 45614 20356 45666
rect 20300 45612 20356 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19852 45106 19908 45108
rect 19852 45054 19854 45106
rect 19854 45054 19906 45106
rect 19906 45054 19908 45106
rect 19852 45052 19908 45054
rect 19964 44828 20020 44884
rect 19292 43820 19348 43876
rect 19516 44268 19572 44324
rect 19628 44044 19684 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19292 43426 19348 43428
rect 19292 43374 19294 43426
rect 19294 43374 19346 43426
rect 19346 43374 19348 43426
rect 19292 43372 19348 43374
rect 19628 43372 19684 43428
rect 19628 42754 19684 42756
rect 19628 42702 19630 42754
rect 19630 42702 19682 42754
rect 19682 42702 19684 42754
rect 19628 42700 19684 42702
rect 19852 43314 19908 43316
rect 19852 43262 19854 43314
rect 19854 43262 19906 43314
rect 19906 43262 19908 43314
rect 19852 43260 19908 43262
rect 20300 42588 20356 42644
rect 19740 42530 19796 42532
rect 19740 42478 19742 42530
rect 19742 42478 19794 42530
rect 19794 42478 19796 42530
rect 19740 42476 19796 42478
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18060 40908 18116 40964
rect 17724 40514 17780 40516
rect 17724 40462 17726 40514
rect 17726 40462 17778 40514
rect 17778 40462 17780 40514
rect 17724 40460 17780 40462
rect 17948 40460 18004 40516
rect 17612 39452 17668 39508
rect 18396 41916 18452 41972
rect 19180 41804 19236 41860
rect 18284 41356 18340 41412
rect 18844 41410 18900 41412
rect 18844 41358 18846 41410
rect 18846 41358 18898 41410
rect 18898 41358 18900 41410
rect 18844 41356 18900 41358
rect 18396 41020 18452 41076
rect 18620 40908 18676 40964
rect 18732 40514 18788 40516
rect 18732 40462 18734 40514
rect 18734 40462 18786 40514
rect 18786 40462 18788 40514
rect 18732 40460 18788 40462
rect 18060 40124 18116 40180
rect 18956 40124 19012 40180
rect 18396 39564 18452 39620
rect 19180 40012 19236 40068
rect 18956 39506 19012 39508
rect 18956 39454 18958 39506
rect 18958 39454 19010 39506
rect 19010 39454 19012 39506
rect 18956 39452 19012 39454
rect 18732 39228 18788 39284
rect 17276 38892 17332 38948
rect 17164 38050 17220 38052
rect 17164 37998 17166 38050
rect 17166 37998 17218 38050
rect 17218 37998 17220 38050
rect 17164 37996 17220 37998
rect 18284 39004 18340 39060
rect 18060 37660 18116 37716
rect 18508 39004 18564 39060
rect 18396 38780 18452 38836
rect 18508 37660 18564 37716
rect 17500 37100 17556 37156
rect 17388 36092 17444 36148
rect 17724 36988 17780 37044
rect 17612 36706 17668 36708
rect 17612 36654 17614 36706
rect 17614 36654 17666 36706
rect 17666 36654 17668 36706
rect 17612 36652 17668 36654
rect 18620 37436 18676 37492
rect 16604 33346 16660 33348
rect 16604 33294 16606 33346
rect 16606 33294 16658 33346
rect 16658 33294 16660 33346
rect 16604 33292 16660 33294
rect 17052 33180 17108 33236
rect 16492 32620 16548 32676
rect 16604 32956 16660 33012
rect 16380 31276 16436 31332
rect 15820 31164 15876 31220
rect 17052 32508 17108 32564
rect 18060 35586 18116 35588
rect 18060 35534 18062 35586
rect 18062 35534 18114 35586
rect 18114 35534 18116 35586
rect 18060 35532 18116 35534
rect 17836 35420 17892 35476
rect 17724 34354 17780 34356
rect 17724 34302 17726 34354
rect 17726 34302 17778 34354
rect 17778 34302 17780 34354
rect 17724 34300 17780 34302
rect 18060 35308 18116 35364
rect 17948 34690 18004 34692
rect 17948 34638 17950 34690
rect 17950 34638 18002 34690
rect 18002 34638 18004 34690
rect 17948 34636 18004 34638
rect 17836 32844 17892 32900
rect 18396 36764 18452 36820
rect 19068 39228 19124 39284
rect 18844 37548 18900 37604
rect 18956 37436 19012 37492
rect 18844 36988 18900 37044
rect 18956 36764 19012 36820
rect 18620 36482 18676 36484
rect 18620 36430 18622 36482
rect 18622 36430 18674 36482
rect 18674 36430 18676 36482
rect 18620 36428 18676 36430
rect 18508 35698 18564 35700
rect 18508 35646 18510 35698
rect 18510 35646 18562 35698
rect 18562 35646 18564 35698
rect 18508 35644 18564 35646
rect 18620 34748 18676 34804
rect 18620 33180 18676 33236
rect 18508 33068 18564 33124
rect 17948 32732 18004 32788
rect 18844 36540 18900 36596
rect 18844 34300 18900 34356
rect 18844 33516 18900 33572
rect 18844 32956 18900 33012
rect 19852 42028 19908 42084
rect 20524 44492 20580 44548
rect 20972 43596 21028 43652
rect 20636 42530 20692 42532
rect 20636 42478 20638 42530
rect 20638 42478 20690 42530
rect 20690 42478 20692 42530
rect 20636 42476 20692 42478
rect 20860 42530 20916 42532
rect 20860 42478 20862 42530
rect 20862 42478 20914 42530
rect 20914 42478 20916 42530
rect 20860 42476 20916 42478
rect 20524 42252 20580 42308
rect 20972 42252 21028 42308
rect 19964 41356 20020 41412
rect 20412 41692 20468 41748
rect 19740 41074 19796 41076
rect 19740 41022 19742 41074
rect 19742 41022 19794 41074
rect 19794 41022 19796 41074
rect 19740 41020 19796 41022
rect 19516 40908 19572 40964
rect 20300 40962 20356 40964
rect 20300 40910 20302 40962
rect 20302 40910 20354 40962
rect 20354 40910 20356 40962
rect 20300 40908 20356 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19852 40402 19908 40404
rect 19852 40350 19854 40402
rect 19854 40350 19906 40402
rect 19906 40350 19908 40402
rect 19852 40348 19908 40350
rect 19516 40012 19572 40068
rect 19404 39900 19460 39956
rect 19964 40124 20020 40180
rect 19964 39730 20020 39732
rect 19964 39678 19966 39730
rect 19966 39678 20018 39730
rect 20018 39678 20020 39730
rect 19964 39676 20020 39678
rect 20300 40124 20356 40180
rect 20972 41580 21028 41636
rect 20748 40684 20804 40740
rect 20524 40348 20580 40404
rect 20636 40236 20692 40292
rect 20524 39618 20580 39620
rect 20524 39566 20526 39618
rect 20526 39566 20578 39618
rect 20578 39566 20580 39618
rect 20524 39564 20580 39566
rect 20412 39340 20468 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19628 38780 19684 38836
rect 19292 38108 19348 38164
rect 19516 37436 19572 37492
rect 19740 38108 19796 38164
rect 19740 37884 19796 37940
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19292 37212 19348 37268
rect 19516 37212 19572 37268
rect 19404 36428 19460 36484
rect 19292 35420 19348 35476
rect 19180 35196 19236 35252
rect 19852 37100 19908 37156
rect 19180 34802 19236 34804
rect 19180 34750 19182 34802
rect 19182 34750 19234 34802
rect 19234 34750 19236 34802
rect 19180 34748 19236 34750
rect 18956 32732 19012 32788
rect 19628 36988 19684 37044
rect 20412 38556 20468 38612
rect 21644 47180 21700 47236
rect 21308 47068 21364 47124
rect 21308 46786 21364 46788
rect 21308 46734 21310 46786
rect 21310 46734 21362 46786
rect 21362 46734 21364 46786
rect 21308 46732 21364 46734
rect 21420 46508 21476 46564
rect 21308 44322 21364 44324
rect 21308 44270 21310 44322
rect 21310 44270 21362 44322
rect 21362 44270 21364 44322
rect 21308 44268 21364 44270
rect 21308 42924 21364 42980
rect 21420 42140 21476 42196
rect 22652 54124 22708 54180
rect 23324 55020 23380 55076
rect 23324 54514 23380 54516
rect 23324 54462 23326 54514
rect 23326 54462 23378 54514
rect 23378 54462 23380 54514
rect 23324 54460 23380 54462
rect 24892 54796 24948 54852
rect 23660 54572 23716 54628
rect 22876 54124 22932 54180
rect 22316 53452 22372 53508
rect 22540 53730 22596 53732
rect 22540 53678 22542 53730
rect 22542 53678 22594 53730
rect 22594 53678 22596 53730
rect 22540 53676 22596 53678
rect 22092 52220 22148 52276
rect 22316 51996 22372 52052
rect 22764 53170 22820 53172
rect 22764 53118 22766 53170
rect 22766 53118 22818 53170
rect 22818 53118 22820 53170
rect 22764 53116 22820 53118
rect 22540 52946 22596 52948
rect 22540 52894 22542 52946
rect 22542 52894 22594 52946
rect 22594 52894 22596 52946
rect 22540 52892 22596 52894
rect 22092 50594 22148 50596
rect 22092 50542 22094 50594
rect 22094 50542 22146 50594
rect 22146 50542 22148 50594
rect 22092 50540 22148 50542
rect 22540 51100 22596 51156
rect 22316 50594 22372 50596
rect 22316 50542 22318 50594
rect 22318 50542 22370 50594
rect 22370 50542 22372 50594
rect 22316 50540 22372 50542
rect 22652 51324 22708 51380
rect 25116 54460 25172 54516
rect 23884 53842 23940 53844
rect 23884 53790 23886 53842
rect 23886 53790 23938 53842
rect 23938 53790 23940 53842
rect 23884 53788 23940 53790
rect 23436 53676 23492 53732
rect 25228 53788 25284 53844
rect 23100 53116 23156 53172
rect 22988 52386 23044 52388
rect 22988 52334 22990 52386
rect 22990 52334 23042 52386
rect 23042 52334 23044 52386
rect 22988 52332 23044 52334
rect 23324 53452 23380 53508
rect 23212 52892 23268 52948
rect 23212 52332 23268 52388
rect 23100 52220 23156 52276
rect 23436 53228 23492 53284
rect 23996 52162 24052 52164
rect 23996 52110 23998 52162
rect 23998 52110 24050 52162
rect 24050 52110 24052 52162
rect 23996 52108 24052 52110
rect 23772 51996 23828 52052
rect 22988 51602 23044 51604
rect 22988 51550 22990 51602
rect 22990 51550 23042 51602
rect 23042 51550 23044 51602
rect 22988 51548 23044 51550
rect 23884 51938 23940 51940
rect 23884 51886 23886 51938
rect 23886 51886 23938 51938
rect 23938 51886 23940 51938
rect 23884 51884 23940 51886
rect 47740 56252 47796 56308
rect 31164 56082 31220 56084
rect 31164 56030 31166 56082
rect 31166 56030 31218 56082
rect 31218 56030 31220 56082
rect 31164 56028 31220 56030
rect 32284 56082 32340 56084
rect 32284 56030 32286 56082
rect 32286 56030 32338 56082
rect 32338 56030 32340 56082
rect 32284 56028 32340 56030
rect 31612 55692 31668 55748
rect 25340 53228 25396 53284
rect 25900 54514 25956 54516
rect 25900 54462 25902 54514
rect 25902 54462 25954 54514
rect 25954 54462 25956 54514
rect 25900 54460 25956 54462
rect 25676 54402 25732 54404
rect 25676 54350 25678 54402
rect 25678 54350 25730 54402
rect 25730 54350 25732 54402
rect 25676 54348 25732 54350
rect 25564 54290 25620 54292
rect 25564 54238 25566 54290
rect 25566 54238 25618 54290
rect 25618 54238 25620 54290
rect 25564 54236 25620 54238
rect 25564 53900 25620 53956
rect 25788 53788 25844 53844
rect 25116 53116 25172 53172
rect 23884 51602 23940 51604
rect 23884 51550 23886 51602
rect 23886 51550 23938 51602
rect 23938 51550 23940 51602
rect 23884 51548 23940 51550
rect 23660 51490 23716 51492
rect 23660 51438 23662 51490
rect 23662 51438 23714 51490
rect 23714 51438 23716 51490
rect 23660 51436 23716 51438
rect 24108 51378 24164 51380
rect 24108 51326 24110 51378
rect 24110 51326 24162 51378
rect 24162 51326 24164 51378
rect 24108 51324 24164 51326
rect 23212 50988 23268 51044
rect 23884 51100 23940 51156
rect 25004 51884 25060 51940
rect 23212 50540 23268 50596
rect 23996 50540 24052 50596
rect 22652 50482 22708 50484
rect 22652 50430 22654 50482
rect 22654 50430 22706 50482
rect 22706 50430 22708 50482
rect 22652 50428 22708 50430
rect 23100 50482 23156 50484
rect 23100 50430 23102 50482
rect 23102 50430 23154 50482
rect 23154 50430 23156 50482
rect 23100 50428 23156 50430
rect 22428 49810 22484 49812
rect 22428 49758 22430 49810
rect 22430 49758 22482 49810
rect 22482 49758 22484 49810
rect 22428 49756 22484 49758
rect 22652 49756 22708 49812
rect 22428 49532 22484 49588
rect 22204 47180 22260 47236
rect 22316 47964 22372 48020
rect 22092 46396 22148 46452
rect 21868 45890 21924 45892
rect 21868 45838 21870 45890
rect 21870 45838 21922 45890
rect 21922 45838 21924 45890
rect 21868 45836 21924 45838
rect 22204 45276 22260 45332
rect 22092 44994 22148 44996
rect 22092 44942 22094 44994
rect 22094 44942 22146 44994
rect 22146 44942 22148 44994
rect 22092 44940 22148 44942
rect 21868 44492 21924 44548
rect 21756 44322 21812 44324
rect 21756 44270 21758 44322
rect 21758 44270 21810 44322
rect 21810 44270 21812 44322
rect 21756 44268 21812 44270
rect 22092 44044 22148 44100
rect 21756 43820 21812 43876
rect 21644 42866 21700 42868
rect 21644 42814 21646 42866
rect 21646 42814 21698 42866
rect 21698 42814 21700 42866
rect 21644 42812 21700 42814
rect 21756 42754 21812 42756
rect 21756 42702 21758 42754
rect 21758 42702 21810 42754
rect 21810 42702 21812 42754
rect 21756 42700 21812 42702
rect 21644 42194 21700 42196
rect 21644 42142 21646 42194
rect 21646 42142 21698 42194
rect 21698 42142 21700 42194
rect 21644 42140 21700 42142
rect 21196 40908 21252 40964
rect 21532 41356 21588 41412
rect 21532 41020 21588 41076
rect 22988 49586 23044 49588
rect 22988 49534 22990 49586
rect 22990 49534 23042 49586
rect 23042 49534 23044 49586
rect 22988 49532 23044 49534
rect 23772 49532 23828 49588
rect 23212 49196 23268 49252
rect 22876 48972 22932 49028
rect 23212 48802 23268 48804
rect 23212 48750 23214 48802
rect 23214 48750 23266 48802
rect 23266 48750 23268 48802
rect 23212 48748 23268 48750
rect 22540 48636 22596 48692
rect 23884 49196 23940 49252
rect 24108 49756 24164 49812
rect 24220 49698 24276 49700
rect 24220 49646 24222 49698
rect 24222 49646 24274 49698
rect 24274 49646 24276 49698
rect 24220 49644 24276 49646
rect 22652 48188 22708 48244
rect 23548 48188 23604 48244
rect 23548 48018 23604 48020
rect 23548 47966 23550 48018
rect 23550 47966 23602 48018
rect 23602 47966 23604 48018
rect 23548 47964 23604 47966
rect 22764 47516 22820 47572
rect 22540 47404 22596 47460
rect 22540 46396 22596 46452
rect 22876 47234 22932 47236
rect 22876 47182 22878 47234
rect 22878 47182 22930 47234
rect 22930 47182 22932 47234
rect 22876 47180 22932 47182
rect 23324 47234 23380 47236
rect 23324 47182 23326 47234
rect 23326 47182 23378 47234
rect 23378 47182 23380 47234
rect 23324 47180 23380 47182
rect 24332 48748 24388 48804
rect 24892 51548 24948 51604
rect 25340 52274 25396 52276
rect 25340 52222 25342 52274
rect 25342 52222 25394 52274
rect 25394 52222 25396 52274
rect 25340 52220 25396 52222
rect 25340 52050 25396 52052
rect 25340 51998 25342 52050
rect 25342 51998 25394 52050
rect 25394 51998 25396 52050
rect 25340 51996 25396 51998
rect 25004 51436 25060 51492
rect 25004 51212 25060 51268
rect 24668 49420 24724 49476
rect 24556 48636 24612 48692
rect 24668 47964 24724 48020
rect 23548 47068 23604 47124
rect 23436 46956 23492 47012
rect 23324 46844 23380 46900
rect 22988 46732 23044 46788
rect 22428 46284 22484 46340
rect 23100 46060 23156 46116
rect 22428 44268 22484 44324
rect 22540 45052 22596 45108
rect 22652 44994 22708 44996
rect 22652 44942 22654 44994
rect 22654 44942 22706 44994
rect 22706 44942 22708 44994
rect 22652 44940 22708 44942
rect 22764 44604 22820 44660
rect 22652 44156 22708 44212
rect 22652 41970 22708 41972
rect 22652 41918 22654 41970
rect 22654 41918 22706 41970
rect 22706 41918 22708 41970
rect 22652 41916 22708 41918
rect 21980 41244 22036 41300
rect 21084 39004 21140 39060
rect 20972 38220 21028 38276
rect 20412 37548 20468 37604
rect 20412 37212 20468 37268
rect 21532 40236 21588 40292
rect 21532 39564 21588 39620
rect 21644 39788 21700 39844
rect 21420 39004 21476 39060
rect 21308 38556 21364 38612
rect 20300 36988 20356 37044
rect 20524 36988 20580 37044
rect 20076 36316 20132 36372
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20300 35868 20356 35924
rect 19964 35026 20020 35028
rect 19964 34974 19966 35026
rect 19966 34974 20018 35026
rect 20018 34974 20020 35026
rect 19964 34972 20020 34974
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20636 34972 20692 35028
rect 20972 35980 21028 36036
rect 22428 41020 22484 41076
rect 22316 40572 22372 40628
rect 22428 40348 22484 40404
rect 23772 46898 23828 46900
rect 23772 46846 23774 46898
rect 23774 46846 23826 46898
rect 23826 46846 23828 46898
rect 23772 46844 23828 46846
rect 23660 46786 23716 46788
rect 23660 46734 23662 46786
rect 23662 46734 23714 46786
rect 23714 46734 23716 46786
rect 23660 46732 23716 46734
rect 23884 46786 23940 46788
rect 23884 46734 23886 46786
rect 23886 46734 23938 46786
rect 23938 46734 23940 46786
rect 23884 46732 23940 46734
rect 23884 46172 23940 46228
rect 24108 47180 24164 47236
rect 24220 47068 24276 47124
rect 23436 46060 23492 46116
rect 23436 44828 23492 44884
rect 23660 44882 23716 44884
rect 23660 44830 23662 44882
rect 23662 44830 23714 44882
rect 23714 44830 23716 44882
rect 23660 44828 23716 44830
rect 23100 44716 23156 44772
rect 23660 44492 23716 44548
rect 23660 44322 23716 44324
rect 23660 44270 23662 44322
rect 23662 44270 23714 44322
rect 23714 44270 23716 44322
rect 23660 44268 23716 44270
rect 23324 44156 23380 44212
rect 22876 42924 22932 42980
rect 23324 43484 23380 43540
rect 23548 44044 23604 44100
rect 22988 43372 23044 43428
rect 22876 42140 22932 42196
rect 23436 42924 23492 42980
rect 24556 46786 24612 46788
rect 24556 46734 24558 46786
rect 24558 46734 24610 46786
rect 24610 46734 24612 46786
rect 24556 46732 24612 46734
rect 24444 46508 24500 46564
rect 24444 45500 24500 45556
rect 24444 45218 24500 45220
rect 24444 45166 24446 45218
rect 24446 45166 24498 45218
rect 24498 45166 24500 45218
rect 24444 45164 24500 45166
rect 24332 45106 24388 45108
rect 24332 45054 24334 45106
rect 24334 45054 24386 45106
rect 24386 45054 24388 45106
rect 24332 45052 24388 45054
rect 24444 44268 24500 44324
rect 24780 47458 24836 47460
rect 24780 47406 24782 47458
rect 24782 47406 24834 47458
rect 24834 47406 24836 47458
rect 24780 47404 24836 47406
rect 23884 43596 23940 43652
rect 22988 42028 23044 42084
rect 23548 42364 23604 42420
rect 23212 41858 23268 41860
rect 23212 41806 23214 41858
rect 23214 41806 23266 41858
rect 23266 41806 23268 41858
rect 23212 41804 23268 41806
rect 22764 40796 22820 40852
rect 22988 40572 23044 40628
rect 22764 39058 22820 39060
rect 22764 39006 22766 39058
rect 22766 39006 22818 39058
rect 22818 39006 22820 39058
rect 22764 39004 22820 39006
rect 21980 37772 22036 37828
rect 21756 37100 21812 37156
rect 21980 36988 22036 37044
rect 21868 36652 21924 36708
rect 21756 36428 21812 36484
rect 21420 35532 21476 35588
rect 21868 35420 21924 35476
rect 20300 34412 20356 34468
rect 19852 34242 19908 34244
rect 19852 34190 19854 34242
rect 19854 34190 19906 34242
rect 19906 34190 19908 34242
rect 19852 34188 19908 34190
rect 19516 33570 19572 33572
rect 19516 33518 19518 33570
rect 19518 33518 19570 33570
rect 19570 33518 19572 33570
rect 19516 33516 19572 33518
rect 17164 31836 17220 31892
rect 16716 31164 16772 31220
rect 15260 29986 15316 29988
rect 15260 29934 15262 29986
rect 15262 29934 15314 29986
rect 15314 29934 15316 29986
rect 15260 29932 15316 29934
rect 18284 31836 18340 31892
rect 18844 31890 18900 31892
rect 18844 31838 18846 31890
rect 18846 31838 18898 31890
rect 18898 31838 18900 31890
rect 18844 31836 18900 31838
rect 19068 31836 19124 31892
rect 19180 33180 19236 33236
rect 18060 31052 18116 31108
rect 17388 30268 17444 30324
rect 16492 29932 16548 29988
rect 18172 30994 18228 30996
rect 18172 30942 18174 30994
rect 18174 30942 18226 30994
rect 18226 30942 18228 30994
rect 18172 30940 18228 30942
rect 17948 30268 18004 30324
rect 17836 30210 17892 30212
rect 17836 30158 17838 30210
rect 17838 30158 17890 30210
rect 17890 30158 17892 30210
rect 17836 30156 17892 30158
rect 23212 39394 23268 39396
rect 23212 39342 23214 39394
rect 23214 39342 23266 39394
rect 23266 39342 23268 39394
rect 23212 39340 23268 39342
rect 23436 38834 23492 38836
rect 23436 38782 23438 38834
rect 23438 38782 23490 38834
rect 23490 38782 23492 38834
rect 23436 38780 23492 38782
rect 22876 38162 22932 38164
rect 22876 38110 22878 38162
rect 22878 38110 22930 38162
rect 22930 38110 22932 38162
rect 22876 38108 22932 38110
rect 22764 37996 22820 38052
rect 23212 37996 23268 38052
rect 23324 38108 23380 38164
rect 22764 37660 22820 37716
rect 22764 36988 22820 37044
rect 22204 34860 22260 34916
rect 22540 34972 22596 35028
rect 20636 34076 20692 34132
rect 20300 33516 20356 33572
rect 20300 33292 20356 33348
rect 20188 33180 20244 33236
rect 19292 33122 19348 33124
rect 19292 33070 19294 33122
rect 19294 33070 19346 33122
rect 19346 33070 19348 33122
rect 19292 33068 19348 33070
rect 19836 32954 19892 32956
rect 19404 32844 19460 32900
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19292 32732 19348 32788
rect 20972 34018 21028 34020
rect 20972 33966 20974 34018
rect 20974 33966 21026 34018
rect 21026 33966 21028 34018
rect 20972 33964 21028 33966
rect 22316 34188 22372 34244
rect 21308 33516 21364 33572
rect 21756 33628 21812 33684
rect 22316 33628 22372 33684
rect 20748 33292 20804 33348
rect 21756 33292 21812 33348
rect 20748 33122 20804 33124
rect 20748 33070 20750 33122
rect 20750 33070 20802 33122
rect 20802 33070 20804 33122
rect 20748 33068 20804 33070
rect 19964 32562 20020 32564
rect 19964 32510 19966 32562
rect 19966 32510 20018 32562
rect 20018 32510 20020 32562
rect 19964 32508 20020 32510
rect 21308 32508 21364 32564
rect 19292 31724 19348 31780
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19180 31164 19236 31220
rect 19740 31218 19796 31220
rect 19740 31166 19742 31218
rect 19742 31166 19794 31218
rect 19794 31166 19796 31218
rect 19740 31164 19796 31166
rect 20300 31218 20356 31220
rect 20300 31166 20302 31218
rect 20302 31166 20354 31218
rect 20354 31166 20356 31218
rect 20300 31164 20356 31166
rect 19628 31106 19684 31108
rect 19628 31054 19630 31106
rect 19630 31054 19682 31106
rect 19682 31054 19684 31106
rect 19628 31052 19684 31054
rect 21532 32732 21588 32788
rect 22204 33068 22260 33124
rect 21756 32060 21812 32116
rect 22428 32786 22484 32788
rect 22428 32734 22430 32786
rect 22430 32734 22482 32786
rect 22482 32734 22484 32786
rect 22428 32732 22484 32734
rect 22652 34130 22708 34132
rect 22652 34078 22654 34130
rect 22654 34078 22706 34130
rect 22706 34078 22708 34130
rect 22652 34076 22708 34078
rect 23660 42642 23716 42644
rect 23660 42590 23662 42642
rect 23662 42590 23714 42642
rect 23714 42590 23716 42642
rect 23660 42588 23716 42590
rect 23660 42028 23716 42084
rect 23772 41692 23828 41748
rect 23996 41356 24052 41412
rect 25228 50876 25284 50932
rect 25340 51324 25396 51380
rect 25900 53506 25956 53508
rect 25900 53454 25902 53506
rect 25902 53454 25954 53506
rect 25954 53454 25956 53506
rect 25900 53452 25956 53454
rect 25564 52444 25620 52500
rect 25676 51602 25732 51604
rect 25676 51550 25678 51602
rect 25678 51550 25730 51602
rect 25730 51550 25732 51602
rect 25676 51548 25732 51550
rect 25788 51378 25844 51380
rect 25788 51326 25790 51378
rect 25790 51326 25842 51378
rect 25842 51326 25844 51378
rect 25788 51324 25844 51326
rect 25564 51100 25620 51156
rect 25564 50594 25620 50596
rect 25564 50542 25566 50594
rect 25566 50542 25618 50594
rect 25618 50542 25620 50594
rect 25564 50540 25620 50542
rect 25228 49644 25284 49700
rect 25228 49420 25284 49476
rect 25900 48188 25956 48244
rect 25116 48076 25172 48132
rect 25564 48076 25620 48132
rect 25228 47292 25284 47348
rect 25004 47068 25060 47124
rect 25340 46898 25396 46900
rect 25340 46846 25342 46898
rect 25342 46846 25394 46898
rect 25394 46846 25396 46898
rect 25340 46844 25396 46846
rect 25228 45778 25284 45780
rect 25228 45726 25230 45778
rect 25230 45726 25282 45778
rect 25282 45726 25284 45778
rect 25228 45724 25284 45726
rect 25004 44828 25060 44884
rect 25340 45276 25396 45332
rect 25452 44828 25508 44884
rect 25340 44322 25396 44324
rect 25340 44270 25342 44322
rect 25342 44270 25394 44322
rect 25394 44270 25396 44322
rect 25340 44268 25396 44270
rect 24220 42700 24276 42756
rect 25676 48018 25732 48020
rect 25676 47966 25678 48018
rect 25678 47966 25730 48018
rect 25730 47966 25732 48018
rect 25676 47964 25732 47966
rect 25676 47628 25732 47684
rect 27468 55074 27524 55076
rect 27468 55022 27470 55074
rect 27470 55022 27522 55074
rect 27522 55022 27524 55074
rect 27468 55020 27524 55022
rect 27916 55074 27972 55076
rect 27916 55022 27918 55074
rect 27918 55022 27970 55074
rect 27970 55022 27972 55074
rect 27916 55020 27972 55022
rect 27132 54514 27188 54516
rect 27132 54462 27134 54514
rect 27134 54462 27186 54514
rect 27186 54462 27188 54514
rect 27132 54460 27188 54462
rect 28588 54796 28644 54852
rect 29372 54796 29428 54852
rect 28028 54684 28084 54740
rect 27244 54236 27300 54292
rect 27804 54012 27860 54068
rect 26124 48524 26180 48580
rect 26124 47404 26180 47460
rect 25900 46844 25956 46900
rect 25788 46396 25844 46452
rect 25676 45836 25732 45892
rect 25788 45388 25844 45444
rect 25676 44828 25732 44884
rect 25228 43538 25284 43540
rect 25228 43486 25230 43538
rect 25230 43486 25282 43538
rect 25282 43486 25284 43538
rect 25228 43484 25284 43486
rect 25564 43426 25620 43428
rect 25564 43374 25566 43426
rect 25566 43374 25618 43426
rect 25618 43374 25620 43426
rect 25564 43372 25620 43374
rect 25452 43314 25508 43316
rect 25452 43262 25454 43314
rect 25454 43262 25506 43314
rect 25506 43262 25508 43314
rect 25452 43260 25508 43262
rect 24668 42754 24724 42756
rect 24668 42702 24670 42754
rect 24670 42702 24722 42754
rect 24722 42702 24724 42754
rect 24668 42700 24724 42702
rect 24892 42700 24948 42756
rect 23660 39116 23716 39172
rect 23660 38834 23716 38836
rect 23660 38782 23662 38834
rect 23662 38782 23714 38834
rect 23714 38782 23716 38834
rect 23660 38780 23716 38782
rect 23548 37826 23604 37828
rect 23548 37774 23550 37826
rect 23550 37774 23602 37826
rect 23602 37774 23604 37826
rect 23548 37772 23604 37774
rect 23548 36482 23604 36484
rect 23548 36430 23550 36482
rect 23550 36430 23602 36482
rect 23602 36430 23604 36482
rect 23548 36428 23604 36430
rect 24108 40460 24164 40516
rect 24108 39730 24164 39732
rect 24108 39678 24110 39730
rect 24110 39678 24162 39730
rect 24162 39678 24164 39730
rect 24108 39676 24164 39678
rect 24220 39340 24276 39396
rect 23996 39004 24052 39060
rect 24108 38946 24164 38948
rect 24108 38894 24110 38946
rect 24110 38894 24162 38946
rect 24162 38894 24164 38946
rect 24108 38892 24164 38894
rect 24108 38108 24164 38164
rect 23772 37436 23828 37492
rect 23660 35980 23716 36036
rect 23548 35922 23604 35924
rect 23548 35870 23550 35922
rect 23550 35870 23602 35922
rect 23602 35870 23604 35922
rect 23548 35868 23604 35870
rect 23436 35644 23492 35700
rect 23436 34860 23492 34916
rect 23212 33852 23268 33908
rect 22876 33740 22932 33796
rect 22652 33346 22708 33348
rect 22652 33294 22654 33346
rect 22654 33294 22706 33346
rect 22706 33294 22708 33346
rect 22652 33292 22708 33294
rect 22876 32674 22932 32676
rect 22876 32622 22878 32674
rect 22878 32622 22930 32674
rect 22930 32622 22932 32674
rect 22876 32620 22932 32622
rect 23100 33292 23156 33348
rect 23324 33292 23380 33348
rect 24108 37884 24164 37940
rect 24332 38332 24388 38388
rect 24556 42252 24612 42308
rect 24780 41970 24836 41972
rect 24780 41918 24782 41970
rect 24782 41918 24834 41970
rect 24834 41918 24836 41970
rect 24780 41916 24836 41918
rect 24556 41746 24612 41748
rect 24556 41694 24558 41746
rect 24558 41694 24610 41746
rect 24610 41694 24612 41746
rect 24556 41692 24612 41694
rect 24444 38556 24500 38612
rect 24444 38108 24500 38164
rect 24556 40460 24612 40516
rect 24332 37772 24388 37828
rect 24332 37548 24388 37604
rect 24332 37266 24388 37268
rect 24332 37214 24334 37266
rect 24334 37214 24386 37266
rect 24386 37214 24388 37266
rect 24332 37212 24388 37214
rect 24444 36876 24500 36932
rect 24668 38722 24724 38724
rect 24668 38670 24670 38722
rect 24670 38670 24722 38722
rect 24722 38670 24724 38722
rect 24668 38668 24724 38670
rect 24668 37826 24724 37828
rect 24668 37774 24670 37826
rect 24670 37774 24722 37826
rect 24722 37774 24724 37826
rect 24668 37772 24724 37774
rect 24892 39506 24948 39508
rect 24892 39454 24894 39506
rect 24894 39454 24946 39506
rect 24946 39454 24948 39506
rect 24892 39452 24948 39454
rect 25004 38162 25060 38164
rect 25004 38110 25006 38162
rect 25006 38110 25058 38162
rect 25058 38110 25060 38162
rect 25004 38108 25060 38110
rect 24892 38050 24948 38052
rect 24892 37998 24894 38050
rect 24894 37998 24946 38050
rect 24946 37998 24948 38050
rect 24892 37996 24948 37998
rect 25676 42588 25732 42644
rect 25228 42364 25284 42420
rect 25564 42252 25620 42308
rect 25452 42028 25508 42084
rect 25228 41356 25284 41412
rect 25340 40514 25396 40516
rect 25340 40462 25342 40514
rect 25342 40462 25394 40514
rect 25394 40462 25396 40514
rect 25340 40460 25396 40462
rect 26124 45276 26180 45332
rect 26908 53506 26964 53508
rect 26908 53454 26910 53506
rect 26910 53454 26962 53506
rect 26962 53454 26964 53506
rect 26908 53452 26964 53454
rect 26796 53228 26852 53284
rect 26460 52444 26516 52500
rect 26460 51378 26516 51380
rect 26460 51326 26462 51378
rect 26462 51326 26514 51378
rect 26514 51326 26516 51378
rect 26460 51324 26516 51326
rect 26460 50482 26516 50484
rect 26460 50430 26462 50482
rect 26462 50430 26514 50482
rect 26514 50430 26516 50482
rect 26460 50428 26516 50430
rect 26684 49644 26740 49700
rect 26460 48412 26516 48468
rect 26460 48242 26516 48244
rect 26460 48190 26462 48242
rect 26462 48190 26514 48242
rect 26514 48190 26516 48242
rect 26460 48188 26516 48190
rect 26348 47852 26404 47908
rect 26236 45052 26292 45108
rect 26908 52162 26964 52164
rect 26908 52110 26910 52162
rect 26910 52110 26962 52162
rect 26962 52110 26964 52162
rect 26908 52108 26964 52110
rect 26908 50428 26964 50484
rect 26908 49420 26964 49476
rect 27692 53506 27748 53508
rect 27692 53454 27694 53506
rect 27694 53454 27746 53506
rect 27746 53454 27748 53506
rect 27692 53452 27748 53454
rect 27356 52220 27412 52276
rect 27244 51938 27300 51940
rect 27244 51886 27246 51938
rect 27246 51886 27298 51938
rect 27298 51886 27300 51938
rect 27244 51884 27300 51886
rect 27132 49868 27188 49924
rect 27132 49196 27188 49252
rect 27244 51100 27300 51156
rect 27020 48972 27076 49028
rect 27132 48412 27188 48468
rect 27356 50540 27412 50596
rect 28476 53842 28532 53844
rect 28476 53790 28478 53842
rect 28478 53790 28530 53842
rect 28530 53790 28532 53842
rect 28476 53788 28532 53790
rect 28252 53452 28308 53508
rect 28140 53228 28196 53284
rect 28812 53228 28868 53284
rect 27692 51996 27748 52052
rect 28588 53004 28644 53060
rect 28252 51436 28308 51492
rect 28364 51324 28420 51380
rect 27580 50706 27636 50708
rect 27580 50654 27582 50706
rect 27582 50654 27634 50706
rect 27634 50654 27636 50706
rect 27580 50652 27636 50654
rect 27804 50540 27860 50596
rect 27356 50316 27412 50372
rect 27356 48636 27412 48692
rect 27468 48972 27524 49028
rect 26908 48130 26964 48132
rect 26908 48078 26910 48130
rect 26910 48078 26962 48130
rect 26962 48078 26964 48130
rect 26908 48076 26964 48078
rect 26012 44268 26068 44324
rect 26684 47068 26740 47124
rect 27356 47570 27412 47572
rect 27356 47518 27358 47570
rect 27358 47518 27410 47570
rect 27410 47518 27412 47570
rect 27356 47516 27412 47518
rect 26796 46732 26852 46788
rect 26460 46396 26516 46452
rect 26572 46284 26628 46340
rect 26796 46396 26852 46452
rect 27468 47292 27524 47348
rect 27580 48412 27636 48468
rect 27580 48188 27636 48244
rect 27020 46620 27076 46676
rect 27356 47180 27412 47236
rect 26684 46060 26740 46116
rect 27020 45890 27076 45892
rect 27020 45838 27022 45890
rect 27022 45838 27074 45890
rect 27074 45838 27076 45890
rect 27020 45836 27076 45838
rect 26572 45388 26628 45444
rect 26684 45330 26740 45332
rect 26684 45278 26686 45330
rect 26686 45278 26738 45330
rect 26738 45278 26740 45330
rect 26684 45276 26740 45278
rect 26348 43484 26404 43540
rect 26796 44994 26852 44996
rect 26796 44942 26798 44994
rect 26798 44942 26850 44994
rect 26850 44942 26852 44994
rect 26796 44940 26852 44942
rect 27244 46674 27300 46676
rect 27244 46622 27246 46674
rect 27246 46622 27298 46674
rect 27298 46622 27300 46674
rect 27244 46620 27300 46622
rect 27132 45164 27188 45220
rect 26908 44604 26964 44660
rect 26908 43596 26964 43652
rect 26684 43260 26740 43316
rect 26124 42476 26180 42532
rect 26012 42364 26068 42420
rect 26572 43036 26628 43092
rect 26012 41970 26068 41972
rect 26012 41918 26014 41970
rect 26014 41918 26066 41970
rect 26066 41918 26068 41970
rect 26012 41916 26068 41918
rect 26572 42028 26628 42084
rect 27468 47068 27524 47124
rect 27692 46508 27748 46564
rect 28252 50652 28308 50708
rect 28140 50482 28196 50484
rect 28140 50430 28142 50482
rect 28142 50430 28194 50482
rect 28194 50430 28196 50482
rect 28140 50428 28196 50430
rect 28476 50428 28532 50484
rect 29484 54572 29540 54628
rect 30156 55132 30212 55188
rect 30828 55186 30884 55188
rect 30828 55134 30830 55186
rect 30830 55134 30882 55186
rect 30882 55134 30884 55186
rect 30828 55132 30884 55134
rect 31500 55132 31556 55188
rect 29708 54460 29764 54516
rect 30156 54402 30212 54404
rect 30156 54350 30158 54402
rect 30158 54350 30210 54402
rect 30210 54350 30212 54402
rect 30156 54348 30212 54350
rect 30044 53900 30100 53956
rect 29260 51436 29316 51492
rect 28812 50316 28868 50372
rect 27916 49644 27972 49700
rect 28028 49810 28084 49812
rect 28028 49758 28030 49810
rect 28030 49758 28082 49810
rect 28082 49758 28084 49810
rect 28028 49756 28084 49758
rect 27916 49196 27972 49252
rect 28588 49698 28644 49700
rect 28588 49646 28590 49698
rect 28590 49646 28642 49698
rect 28642 49646 28644 49698
rect 28588 49644 28644 49646
rect 28028 48972 28084 49028
rect 28812 49084 28868 49140
rect 29148 50594 29204 50596
rect 29148 50542 29150 50594
rect 29150 50542 29202 50594
rect 29202 50542 29204 50594
rect 29148 50540 29204 50542
rect 29708 50370 29764 50372
rect 29708 50318 29710 50370
rect 29710 50318 29762 50370
rect 29762 50318 29764 50370
rect 29708 50316 29764 50318
rect 30380 52668 30436 52724
rect 30156 52556 30212 52612
rect 30156 51324 30212 51380
rect 30604 55020 30660 55076
rect 30940 53788 30996 53844
rect 30828 53170 30884 53172
rect 30828 53118 30830 53170
rect 30830 53118 30882 53170
rect 30882 53118 30884 53170
rect 30828 53116 30884 53118
rect 30940 52834 30996 52836
rect 30940 52782 30942 52834
rect 30942 52782 30994 52834
rect 30994 52782 30996 52834
rect 30940 52780 30996 52782
rect 31164 52668 31220 52724
rect 30828 51996 30884 52052
rect 30044 50540 30100 50596
rect 30268 50316 30324 50372
rect 31276 52050 31332 52052
rect 31276 51998 31278 52050
rect 31278 51998 31330 52050
rect 31330 51998 31332 52050
rect 31276 51996 31332 51998
rect 31164 51660 31220 51716
rect 30940 51436 30996 51492
rect 30828 51378 30884 51380
rect 30828 51326 30830 51378
rect 30830 51326 30882 51378
rect 30882 51326 30884 51378
rect 30828 51324 30884 51326
rect 30716 51212 30772 51268
rect 30492 50316 30548 50372
rect 30044 49922 30100 49924
rect 30044 49870 30046 49922
rect 30046 49870 30098 49922
rect 30098 49870 30100 49922
rect 30044 49868 30100 49870
rect 30268 49810 30324 49812
rect 30268 49758 30270 49810
rect 30270 49758 30322 49810
rect 30322 49758 30324 49810
rect 30268 49756 30324 49758
rect 29708 49644 29764 49700
rect 28588 48802 28644 48804
rect 28588 48750 28590 48802
rect 28590 48750 28642 48802
rect 28642 48750 28644 48802
rect 28588 48748 28644 48750
rect 29148 49420 29204 49476
rect 28028 48188 28084 48244
rect 28364 48188 28420 48244
rect 28140 47458 28196 47460
rect 28140 47406 28142 47458
rect 28142 47406 28194 47458
rect 28194 47406 28196 47458
rect 28140 47404 28196 47406
rect 28252 47346 28308 47348
rect 28252 47294 28254 47346
rect 28254 47294 28306 47346
rect 28306 47294 28308 47346
rect 28252 47292 28308 47294
rect 28364 47068 28420 47124
rect 28028 46956 28084 47012
rect 27916 46284 27972 46340
rect 27804 46172 27860 46228
rect 28028 46172 28084 46228
rect 27692 45948 27748 46004
rect 28364 45890 28420 45892
rect 28364 45838 28366 45890
rect 28366 45838 28418 45890
rect 28418 45838 28420 45890
rect 28364 45836 28420 45838
rect 28140 45666 28196 45668
rect 28140 45614 28142 45666
rect 28142 45614 28194 45666
rect 28194 45614 28196 45666
rect 28140 45612 28196 45614
rect 27468 45106 27524 45108
rect 27468 45054 27470 45106
rect 27470 45054 27522 45106
rect 27522 45054 27524 45106
rect 27468 45052 27524 45054
rect 27580 43538 27636 43540
rect 27580 43486 27582 43538
rect 27582 43486 27634 43538
rect 27634 43486 27636 43538
rect 27580 43484 27636 43486
rect 27580 43260 27636 43316
rect 26796 42028 26852 42084
rect 26348 41804 26404 41860
rect 25788 40012 25844 40068
rect 25228 39340 25284 39396
rect 25340 38556 25396 38612
rect 26124 40796 26180 40852
rect 26236 40684 26292 40740
rect 26684 41804 26740 41860
rect 26012 39004 26068 39060
rect 26236 39116 26292 39172
rect 26124 38892 26180 38948
rect 26348 39004 26404 39060
rect 26124 38668 26180 38724
rect 26572 41356 26628 41412
rect 26796 40514 26852 40516
rect 26796 40462 26798 40514
rect 26798 40462 26850 40514
rect 26850 40462 26852 40514
rect 26796 40460 26852 40462
rect 25676 38332 25732 38388
rect 24780 37660 24836 37716
rect 25116 37548 25172 37604
rect 25340 38050 25396 38052
rect 25340 37998 25342 38050
rect 25342 37998 25394 38050
rect 25394 37998 25396 38050
rect 25340 37996 25396 37998
rect 25116 36706 25172 36708
rect 25116 36654 25118 36706
rect 25118 36654 25170 36706
rect 25170 36654 25172 36706
rect 25116 36652 25172 36654
rect 24108 35532 24164 35588
rect 24220 35980 24276 36036
rect 23772 34188 23828 34244
rect 23436 33628 23492 33684
rect 23884 33516 23940 33572
rect 23212 32956 23268 33012
rect 23324 33068 23380 33124
rect 23660 33122 23716 33124
rect 23660 33070 23662 33122
rect 23662 33070 23714 33122
rect 23714 33070 23716 33122
rect 23660 33068 23716 33070
rect 25340 36540 25396 36596
rect 24444 36428 24500 36484
rect 25564 37436 25620 37492
rect 24556 36316 24612 36372
rect 25564 36876 25620 36932
rect 24444 35922 24500 35924
rect 24444 35870 24446 35922
rect 24446 35870 24498 35922
rect 24498 35870 24500 35922
rect 24444 35868 24500 35870
rect 24668 35532 24724 35588
rect 25116 35980 25172 36036
rect 24668 34524 24724 34580
rect 24444 34242 24500 34244
rect 24444 34190 24446 34242
rect 24446 34190 24498 34242
rect 24498 34190 24500 34242
rect 24444 34188 24500 34190
rect 24780 34076 24836 34132
rect 24668 33516 24724 33572
rect 24220 33346 24276 33348
rect 24220 33294 24222 33346
rect 24222 33294 24274 33346
rect 24274 33294 24276 33346
rect 24220 33292 24276 33294
rect 24108 32732 24164 32788
rect 24668 32674 24724 32676
rect 24668 32622 24670 32674
rect 24670 32622 24722 32674
rect 24722 32622 24724 32674
rect 24668 32620 24724 32622
rect 24892 33740 24948 33796
rect 24108 32396 24164 32452
rect 23996 31890 24052 31892
rect 23996 31838 23998 31890
rect 23998 31838 24050 31890
rect 24050 31838 24052 31890
rect 23996 31836 24052 31838
rect 23660 31612 23716 31668
rect 20972 30882 21028 30884
rect 20972 30830 20974 30882
rect 20974 30830 21026 30882
rect 21026 30830 21028 30882
rect 20972 30828 21028 30830
rect 16044 28028 16100 28084
rect 16044 27356 16100 27412
rect 15036 27132 15092 27188
rect 13468 26684 13524 26740
rect 14028 26460 14084 26516
rect 12348 25676 12404 25732
rect 14476 26012 14532 26068
rect 12236 24556 12292 24612
rect 9100 23714 9156 23716
rect 9100 23662 9102 23714
rect 9102 23662 9154 23714
rect 9154 23662 9156 23714
rect 9100 23660 9156 23662
rect 10668 24220 10724 24276
rect 9548 23324 9604 23380
rect 10108 23884 10164 23940
rect 8876 23212 8932 23268
rect 8316 23154 8372 23156
rect 8316 23102 8318 23154
rect 8318 23102 8370 23154
rect 8370 23102 8372 23154
rect 8316 23100 8372 23102
rect 8428 22146 8484 22148
rect 8428 22094 8430 22146
rect 8430 22094 8482 22146
rect 8482 22094 8484 22146
rect 8428 22092 8484 22094
rect 7980 21756 8036 21812
rect 7868 20748 7924 20804
rect 7644 19794 7700 19796
rect 7644 19742 7646 19794
rect 7646 19742 7698 19794
rect 7698 19742 7700 19794
rect 7644 19740 7700 19742
rect 7420 19122 7476 19124
rect 7420 19070 7422 19122
rect 7422 19070 7474 19122
rect 7474 19070 7476 19122
rect 7420 19068 7476 19070
rect 7868 18674 7924 18676
rect 7868 18622 7870 18674
rect 7870 18622 7922 18674
rect 7922 18622 7924 18674
rect 7868 18620 7924 18622
rect 6972 18450 7028 18452
rect 6972 18398 6974 18450
rect 6974 18398 7026 18450
rect 7026 18398 7028 18450
rect 6972 18396 7028 18398
rect 7196 18450 7252 18452
rect 7196 18398 7198 18450
rect 7198 18398 7250 18450
rect 7250 18398 7252 18450
rect 7196 18396 7252 18398
rect 6972 16882 7028 16884
rect 6972 16830 6974 16882
rect 6974 16830 7026 16882
rect 7026 16830 7028 16882
rect 6972 16828 7028 16830
rect 7308 16716 7364 16772
rect 7532 17612 7588 17668
rect 6972 15986 7028 15988
rect 6972 15934 6974 15986
rect 6974 15934 7026 15986
rect 7026 15934 7028 15986
rect 6972 15932 7028 15934
rect 7644 16994 7700 16996
rect 7644 16942 7646 16994
rect 7646 16942 7698 16994
rect 7698 16942 7700 16994
rect 7644 16940 7700 16942
rect 7084 15260 7140 15316
rect 6748 14588 6804 14644
rect 6860 14812 6916 14868
rect 6524 13634 6580 13636
rect 6524 13582 6526 13634
rect 6526 13582 6578 13634
rect 6578 13582 6580 13634
rect 6524 13580 6580 13582
rect 6300 12962 6356 12964
rect 6300 12910 6302 12962
rect 6302 12910 6354 12962
rect 6354 12910 6356 12962
rect 6300 12908 6356 12910
rect 6748 13074 6804 13076
rect 6748 13022 6750 13074
rect 6750 13022 6802 13074
rect 6802 13022 6804 13074
rect 6748 13020 6804 13022
rect 6636 12908 6692 12964
rect 6972 14028 7028 14084
rect 6636 10892 6692 10948
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 6076 9996 6132 10052
rect 5964 9938 6020 9940
rect 5964 9886 5966 9938
rect 5966 9886 6018 9938
rect 6018 9886 6020 9938
rect 5964 9884 6020 9886
rect 3276 9548 3332 9604
rect 6524 10610 6580 10612
rect 6524 10558 6526 10610
rect 6526 10558 6578 10610
rect 6578 10558 6580 10610
rect 6524 10556 6580 10558
rect 6188 9212 6244 9268
rect 1708 8764 1764 8820
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 6412 8428 6468 8484
rect 6300 8370 6356 8372
rect 6300 8318 6302 8370
rect 6302 8318 6354 8370
rect 6354 8318 6356 8370
rect 6300 8316 6356 8318
rect 6524 8204 6580 8260
rect 6860 12066 6916 12068
rect 6860 12014 6862 12066
rect 6862 12014 6914 12066
rect 6914 12014 6916 12066
rect 6860 12012 6916 12014
rect 7196 13692 7252 13748
rect 7196 13522 7252 13524
rect 7196 13470 7198 13522
rect 7198 13470 7250 13522
rect 7250 13470 7252 13522
rect 7196 13468 7252 13470
rect 7084 13356 7140 13412
rect 7084 12962 7140 12964
rect 7084 12910 7086 12962
rect 7086 12910 7138 12962
rect 7138 12910 7140 12962
rect 7084 12908 7140 12910
rect 7756 15372 7812 15428
rect 7644 14754 7700 14756
rect 7644 14702 7646 14754
rect 7646 14702 7698 14754
rect 7698 14702 7700 14754
rect 7644 14700 7700 14702
rect 8204 20188 8260 20244
rect 8204 18620 8260 18676
rect 7980 17612 8036 17668
rect 7980 17442 8036 17444
rect 7980 17390 7982 17442
rect 7982 17390 8034 17442
rect 8034 17390 8036 17442
rect 7980 17388 8036 17390
rect 8988 22316 9044 22372
rect 9324 23100 9380 23156
rect 10556 23154 10612 23156
rect 10556 23102 10558 23154
rect 10558 23102 10610 23154
rect 10610 23102 10612 23154
rect 10556 23100 10612 23102
rect 9660 22370 9716 22372
rect 9660 22318 9662 22370
rect 9662 22318 9714 22370
rect 9714 22318 9716 22370
rect 9660 22316 9716 22318
rect 9772 22258 9828 22260
rect 9772 22206 9774 22258
rect 9774 22206 9826 22258
rect 9826 22206 9828 22258
rect 9772 22204 9828 22206
rect 8876 20524 8932 20580
rect 9772 20524 9828 20580
rect 8652 20130 8708 20132
rect 8652 20078 8654 20130
rect 8654 20078 8706 20130
rect 8706 20078 8708 20130
rect 8652 20076 8708 20078
rect 8652 19010 8708 19012
rect 8652 18958 8654 19010
rect 8654 18958 8706 19010
rect 8706 18958 8708 19010
rect 8652 18956 8708 18958
rect 8764 18396 8820 18452
rect 8428 17052 8484 17108
rect 8316 16940 8372 16996
rect 8428 16716 8484 16772
rect 8204 16322 8260 16324
rect 8204 16270 8206 16322
rect 8206 16270 8258 16322
rect 8258 16270 8260 16322
rect 8204 16268 8260 16270
rect 8428 15148 8484 15204
rect 8876 17442 8932 17444
rect 8876 17390 8878 17442
rect 8878 17390 8930 17442
rect 8930 17390 8932 17442
rect 8876 17388 8932 17390
rect 9212 18956 9268 19012
rect 9660 18956 9716 19012
rect 9100 18844 9156 18900
rect 9548 18284 9604 18340
rect 9660 18060 9716 18116
rect 7980 15036 8036 15092
rect 8204 15036 8260 15092
rect 7868 14812 7924 14868
rect 8316 14924 8372 14980
rect 8204 14028 8260 14084
rect 8092 13692 8148 13748
rect 7532 13356 7588 13412
rect 7420 12850 7476 12852
rect 7420 12798 7422 12850
rect 7422 12798 7474 12850
rect 7474 12798 7476 12850
rect 7420 12796 7476 12798
rect 6972 10892 7028 10948
rect 7084 10834 7140 10836
rect 7084 10782 7086 10834
rect 7086 10782 7138 10834
rect 7138 10782 7140 10834
rect 7084 10780 7140 10782
rect 7644 13580 7700 13636
rect 7532 11506 7588 11508
rect 7532 11454 7534 11506
rect 7534 11454 7586 11506
rect 7586 11454 7588 11506
rect 7532 11452 7588 11454
rect 7308 10892 7364 10948
rect 7756 10610 7812 10612
rect 7756 10558 7758 10610
rect 7758 10558 7810 10610
rect 7810 10558 7812 10610
rect 7756 10556 7812 10558
rect 6860 9436 6916 9492
rect 6860 9266 6916 9268
rect 6860 9214 6862 9266
rect 6862 9214 6914 9266
rect 6914 9214 6916 9266
rect 6860 9212 6916 9214
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 6748 6860 6804 6916
rect 7756 9826 7812 9828
rect 7756 9774 7758 9826
rect 7758 9774 7810 9826
rect 7810 9774 7812 9826
rect 7756 9772 7812 9774
rect 8540 13916 8596 13972
rect 8204 13580 8260 13636
rect 8428 12796 8484 12852
rect 8540 13468 8596 13524
rect 8988 16994 9044 16996
rect 8988 16942 8990 16994
rect 8990 16942 9042 16994
rect 9042 16942 9044 16994
rect 8988 16940 9044 16942
rect 9324 16828 9380 16884
rect 11228 23938 11284 23940
rect 11228 23886 11230 23938
rect 11230 23886 11282 23938
rect 11282 23886 11284 23938
rect 11228 23884 11284 23886
rect 11676 23436 11732 23492
rect 10892 22482 10948 22484
rect 10892 22430 10894 22482
rect 10894 22430 10946 22482
rect 10946 22430 10948 22482
rect 10892 22428 10948 22430
rect 10220 22092 10276 22148
rect 10780 22092 10836 22148
rect 10668 20578 10724 20580
rect 10668 20526 10670 20578
rect 10670 20526 10722 20578
rect 10722 20526 10724 20578
rect 10668 20524 10724 20526
rect 9996 20076 10052 20132
rect 10108 19234 10164 19236
rect 10108 19182 10110 19234
rect 10110 19182 10162 19234
rect 10162 19182 10164 19234
rect 10108 19180 10164 19182
rect 9884 18396 9940 18452
rect 9884 17106 9940 17108
rect 9884 17054 9886 17106
rect 9886 17054 9938 17106
rect 9938 17054 9940 17106
rect 9884 17052 9940 17054
rect 9100 14700 9156 14756
rect 9212 14530 9268 14532
rect 9212 14478 9214 14530
rect 9214 14478 9266 14530
rect 9266 14478 9268 14530
rect 9212 14476 9268 14478
rect 8876 13356 8932 13412
rect 7980 12178 8036 12180
rect 7980 12126 7982 12178
rect 7982 12126 8034 12178
rect 8034 12126 8036 12178
rect 7980 12124 8036 12126
rect 8092 10892 8148 10948
rect 7980 10556 8036 10612
rect 7308 7868 7364 7924
rect 7420 8428 7476 8484
rect 7308 6802 7364 6804
rect 7308 6750 7310 6802
rect 7310 6750 7362 6802
rect 7362 6750 7364 6802
rect 7308 6748 7364 6750
rect 7196 5852 7252 5908
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 7756 9212 7812 9268
rect 8428 12460 8484 12516
rect 8316 11954 8372 11956
rect 8316 11902 8318 11954
rect 8318 11902 8370 11954
rect 8370 11902 8372 11954
rect 8316 11900 8372 11902
rect 9100 12402 9156 12404
rect 9100 12350 9102 12402
rect 9102 12350 9154 12402
rect 9154 12350 9156 12402
rect 9100 12348 9156 12350
rect 8988 11788 9044 11844
rect 8540 10780 8596 10836
rect 8764 11506 8820 11508
rect 8764 11454 8766 11506
rect 8766 11454 8818 11506
rect 8818 11454 8820 11506
rect 8764 11452 8820 11454
rect 9324 11170 9380 11172
rect 9324 11118 9326 11170
rect 9326 11118 9378 11170
rect 9378 11118 9380 11170
rect 9324 11116 9380 11118
rect 8316 9154 8372 9156
rect 8316 9102 8318 9154
rect 8318 9102 8370 9154
rect 8370 9102 8372 9154
rect 8316 9100 8372 9102
rect 7644 8316 7700 8372
rect 7644 7196 7700 7252
rect 7756 6972 7812 7028
rect 7756 6188 7812 6244
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 7756 3276 7812 3332
rect 7980 8316 8036 8372
rect 8428 8258 8484 8260
rect 8428 8206 8430 8258
rect 8430 8206 8482 8258
rect 8482 8206 8484 8258
rect 8428 8204 8484 8206
rect 7980 6802 8036 6804
rect 7980 6750 7982 6802
rect 7982 6750 8034 6802
rect 8034 6750 8036 6802
rect 7980 6748 8036 6750
rect 10668 19740 10724 19796
rect 10780 18732 10836 18788
rect 10556 18338 10612 18340
rect 10556 18286 10558 18338
rect 10558 18286 10610 18338
rect 10610 18286 10612 18338
rect 10556 18284 10612 18286
rect 10444 16828 10500 16884
rect 10108 16604 10164 16660
rect 10332 16492 10388 16548
rect 9548 15426 9604 15428
rect 9548 15374 9550 15426
rect 9550 15374 9602 15426
rect 9602 15374 9604 15426
rect 9548 15372 9604 15374
rect 9548 14588 9604 14644
rect 10444 15708 10500 15764
rect 10108 15426 10164 15428
rect 10108 15374 10110 15426
rect 10110 15374 10162 15426
rect 10162 15374 10164 15426
rect 10108 15372 10164 15374
rect 9996 15036 10052 15092
rect 10108 14700 10164 14756
rect 9772 14418 9828 14420
rect 9772 14366 9774 14418
rect 9774 14366 9826 14418
rect 9826 14366 9828 14418
rect 9772 14364 9828 14366
rect 9884 14306 9940 14308
rect 9884 14254 9886 14306
rect 9886 14254 9938 14306
rect 9938 14254 9940 14306
rect 9884 14252 9940 14254
rect 9772 13746 9828 13748
rect 9772 13694 9774 13746
rect 9774 13694 9826 13746
rect 9826 13694 9828 13746
rect 9772 13692 9828 13694
rect 9660 12850 9716 12852
rect 9660 12798 9662 12850
rect 9662 12798 9714 12850
rect 9714 12798 9716 12850
rect 9660 12796 9716 12798
rect 10332 14476 10388 14532
rect 10444 14418 10500 14420
rect 10444 14366 10446 14418
rect 10446 14366 10498 14418
rect 10498 14366 10500 14418
rect 10444 14364 10500 14366
rect 10220 14140 10276 14196
rect 10444 13692 10500 13748
rect 10108 12850 10164 12852
rect 10108 12798 10110 12850
rect 10110 12798 10162 12850
rect 10162 12798 10164 12850
rect 10108 12796 10164 12798
rect 10332 11788 10388 11844
rect 10108 11506 10164 11508
rect 10108 11454 10110 11506
rect 10110 11454 10162 11506
rect 10162 11454 10164 11506
rect 10108 11452 10164 11454
rect 10332 11340 10388 11396
rect 9436 9996 9492 10052
rect 9660 11004 9716 11060
rect 8652 8652 8708 8708
rect 8876 9772 8932 9828
rect 9100 9436 9156 9492
rect 9436 9212 9492 9268
rect 9100 8316 9156 8372
rect 8204 6914 8260 6916
rect 8204 6862 8206 6914
rect 8206 6862 8258 6914
rect 8258 6862 8260 6914
rect 8204 6860 8260 6862
rect 10108 10834 10164 10836
rect 10108 10782 10110 10834
rect 10110 10782 10162 10834
rect 10162 10782 10164 10834
rect 10108 10780 10164 10782
rect 9884 9938 9940 9940
rect 9884 9886 9886 9938
rect 9886 9886 9938 9938
rect 9938 9886 9940 9938
rect 9884 9884 9940 9886
rect 9884 9660 9940 9716
rect 9772 8540 9828 8596
rect 10668 17666 10724 17668
rect 10668 17614 10670 17666
rect 10670 17614 10722 17666
rect 10722 17614 10724 17666
rect 10668 17612 10724 17614
rect 10780 16268 10836 16324
rect 11228 22092 11284 22148
rect 11900 23324 11956 23380
rect 11116 21868 11172 21924
rect 11340 21420 11396 21476
rect 11004 20636 11060 20692
rect 11004 19740 11060 19796
rect 11564 22370 11620 22372
rect 11564 22318 11566 22370
rect 11566 22318 11618 22370
rect 11618 22318 11620 22370
rect 11564 22316 11620 22318
rect 11788 22092 11844 22148
rect 11564 20690 11620 20692
rect 11564 20638 11566 20690
rect 11566 20638 11618 20690
rect 11618 20638 11620 20690
rect 11564 20636 11620 20638
rect 11116 18396 11172 18452
rect 11564 18956 11620 19012
rect 11340 18732 11396 18788
rect 11228 15932 11284 15988
rect 11116 15820 11172 15876
rect 12012 23266 12068 23268
rect 12012 23214 12014 23266
rect 12014 23214 12066 23266
rect 12066 23214 12068 23266
rect 12012 23212 12068 23214
rect 12572 23884 12628 23940
rect 11900 21868 11956 21924
rect 12012 20188 12068 20244
rect 11900 19906 11956 19908
rect 11900 19854 11902 19906
rect 11902 19854 11954 19906
rect 11954 19854 11956 19906
rect 11900 19852 11956 19854
rect 11676 18396 11732 18452
rect 13916 24610 13972 24612
rect 13916 24558 13918 24610
rect 13918 24558 13970 24610
rect 13970 24558 13972 24610
rect 13916 24556 13972 24558
rect 14140 24722 14196 24724
rect 14140 24670 14142 24722
rect 14142 24670 14194 24722
rect 14194 24670 14196 24722
rect 14140 24668 14196 24670
rect 14364 23938 14420 23940
rect 14364 23886 14366 23938
rect 14366 23886 14418 23938
rect 14418 23886 14420 23938
rect 14364 23884 14420 23886
rect 12796 23324 12852 23380
rect 13580 23324 13636 23380
rect 12684 23212 12740 23268
rect 12348 22092 12404 22148
rect 12908 22988 12964 23044
rect 12460 20914 12516 20916
rect 12460 20862 12462 20914
rect 12462 20862 12514 20914
rect 12514 20862 12516 20914
rect 12460 20860 12516 20862
rect 12348 20130 12404 20132
rect 12348 20078 12350 20130
rect 12350 20078 12402 20130
rect 12402 20078 12404 20130
rect 12348 20076 12404 20078
rect 12348 18620 12404 18676
rect 12348 18284 12404 18340
rect 11676 18060 11732 18116
rect 10668 14700 10724 14756
rect 10668 14140 10724 14196
rect 10668 13746 10724 13748
rect 10668 13694 10670 13746
rect 10670 13694 10722 13746
rect 10722 13694 10724 13746
rect 10668 13692 10724 13694
rect 11900 17778 11956 17780
rect 11900 17726 11902 17778
rect 11902 17726 11954 17778
rect 11954 17726 11956 17778
rect 11900 17724 11956 17726
rect 11900 17052 11956 17108
rect 12012 16994 12068 16996
rect 12012 16942 12014 16994
rect 12014 16942 12066 16994
rect 12066 16942 12068 16994
rect 12012 16940 12068 16942
rect 12012 16210 12068 16212
rect 12012 16158 12014 16210
rect 12014 16158 12066 16210
rect 12066 16158 12068 16210
rect 12012 16156 12068 16158
rect 11340 14812 11396 14868
rect 11228 14364 11284 14420
rect 11676 15932 11732 15988
rect 11116 12572 11172 12628
rect 10892 12236 10948 12292
rect 11116 12124 11172 12180
rect 10892 11676 10948 11732
rect 11116 11394 11172 11396
rect 11116 11342 11118 11394
rect 11118 11342 11170 11394
rect 11170 11342 11172 11394
rect 11116 11340 11172 11342
rect 10668 11282 10724 11284
rect 10668 11230 10670 11282
rect 10670 11230 10722 11282
rect 10722 11230 10724 11282
rect 10668 11228 10724 11230
rect 10556 9826 10612 9828
rect 10556 9774 10558 9826
rect 10558 9774 10610 9826
rect 10610 9774 10612 9826
rect 10556 9772 10612 9774
rect 10556 8818 10612 8820
rect 10556 8766 10558 8818
rect 10558 8766 10610 8818
rect 10610 8766 10612 8818
rect 10556 8764 10612 8766
rect 9884 8428 9940 8484
rect 9772 8204 9828 8260
rect 9884 7868 9940 7924
rect 8988 6466 9044 6468
rect 8988 6414 8990 6466
rect 8990 6414 9042 6466
rect 9042 6414 9044 6466
rect 8988 6412 9044 6414
rect 9548 6748 9604 6804
rect 9884 6578 9940 6580
rect 9884 6526 9886 6578
rect 9886 6526 9938 6578
rect 9938 6526 9940 6578
rect 9884 6524 9940 6526
rect 9436 5964 9492 6020
rect 8540 5068 8596 5124
rect 9212 5234 9268 5236
rect 9212 5182 9214 5234
rect 9214 5182 9266 5234
rect 9266 5182 9268 5234
rect 9212 5180 9268 5182
rect 9660 6412 9716 6468
rect 9772 6130 9828 6132
rect 9772 6078 9774 6130
rect 9774 6078 9826 6130
rect 9826 6078 9828 6130
rect 9772 6076 9828 6078
rect 11004 9548 11060 9604
rect 11004 8652 11060 8708
rect 10332 7196 10388 7252
rect 10220 5906 10276 5908
rect 10220 5854 10222 5906
rect 10222 5854 10274 5906
rect 10274 5854 10276 5906
rect 10220 5852 10276 5854
rect 10108 5740 10164 5796
rect 10108 4508 10164 4564
rect 10780 7362 10836 7364
rect 10780 7310 10782 7362
rect 10782 7310 10834 7362
rect 10834 7310 10836 7362
rect 10780 7308 10836 7310
rect 10668 6636 10724 6692
rect 10668 5516 10724 5572
rect 10444 4396 10500 4452
rect 10668 4562 10724 4564
rect 10668 4510 10670 4562
rect 10670 4510 10722 4562
rect 10722 4510 10724 4562
rect 10668 4508 10724 4510
rect 10668 3388 10724 3444
rect 11452 13746 11508 13748
rect 11452 13694 11454 13746
rect 11454 13694 11506 13746
rect 11506 13694 11508 13746
rect 11452 13692 11508 13694
rect 11564 13132 11620 13188
rect 11452 12572 11508 12628
rect 11564 12012 11620 12068
rect 12348 16940 12404 16996
rect 12460 16716 12516 16772
rect 11788 15426 11844 15428
rect 11788 15374 11790 15426
rect 11790 15374 11842 15426
rect 11842 15374 11844 15426
rect 11788 15372 11844 15374
rect 11788 15036 11844 15092
rect 11900 14140 11956 14196
rect 12012 13020 12068 13076
rect 11676 11282 11732 11284
rect 11676 11230 11678 11282
rect 11678 11230 11730 11282
rect 11730 11230 11732 11282
rect 11676 11228 11732 11230
rect 11564 10892 11620 10948
rect 11340 9772 11396 9828
rect 11452 9996 11508 10052
rect 11228 9212 11284 9268
rect 11228 8258 11284 8260
rect 11228 8206 11230 8258
rect 11230 8206 11282 8258
rect 11282 8206 11284 8258
rect 11228 8204 11284 8206
rect 11340 7644 11396 7700
rect 11116 6690 11172 6692
rect 11116 6638 11118 6690
rect 11118 6638 11170 6690
rect 11170 6638 11172 6690
rect 11116 6636 11172 6638
rect 11340 6300 11396 6356
rect 11452 7084 11508 7140
rect 11676 10668 11732 10724
rect 11788 10444 11844 10500
rect 13020 22428 13076 22484
rect 12908 22146 12964 22148
rect 12908 22094 12910 22146
rect 12910 22094 12962 22146
rect 12962 22094 12964 22146
rect 12908 22092 12964 22094
rect 13468 22092 13524 22148
rect 13244 21474 13300 21476
rect 13244 21422 13246 21474
rect 13246 21422 13298 21474
rect 13298 21422 13300 21474
rect 13244 21420 13300 21422
rect 13468 20860 13524 20916
rect 12908 19010 12964 19012
rect 12908 18958 12910 19010
rect 12910 18958 12962 19010
rect 12962 18958 12964 19010
rect 12908 18956 12964 18958
rect 12908 18732 12964 18788
rect 12796 18508 12852 18564
rect 13020 17500 13076 17556
rect 12908 16380 12964 16436
rect 12796 15036 12852 15092
rect 12684 14140 12740 14196
rect 13580 20412 13636 20468
rect 13916 23100 13972 23156
rect 13916 22316 13972 22372
rect 14252 21756 14308 21812
rect 13804 20860 13860 20916
rect 14028 20300 14084 20356
rect 13692 18620 13748 18676
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 13580 17724 13636 17780
rect 13468 16716 13524 16772
rect 13468 16492 13524 16548
rect 13356 16156 13412 16212
rect 12796 13804 12852 13860
rect 13020 13916 13076 13972
rect 12348 12738 12404 12740
rect 12348 12686 12350 12738
rect 12350 12686 12402 12738
rect 12402 12686 12404 12738
rect 12348 12684 12404 12686
rect 12236 12572 12292 12628
rect 12236 12348 12292 12404
rect 12572 12348 12628 12404
rect 12124 12236 12180 12292
rect 12012 12012 12068 12068
rect 12012 11788 12068 11844
rect 12124 10556 12180 10612
rect 11900 9042 11956 9044
rect 11900 8990 11902 9042
rect 11902 8990 11954 9042
rect 11954 8990 11956 9042
rect 11900 8988 11956 8990
rect 11788 7868 11844 7924
rect 11676 6972 11732 7028
rect 11452 6748 11508 6804
rect 10892 4508 10948 4564
rect 11676 6748 11732 6804
rect 12236 9826 12292 9828
rect 12236 9774 12238 9826
rect 12238 9774 12290 9826
rect 12290 9774 12292 9826
rect 12236 9772 12292 9774
rect 12684 12178 12740 12180
rect 12684 12126 12686 12178
rect 12686 12126 12738 12178
rect 12738 12126 12740 12178
rect 12684 12124 12740 12126
rect 12572 11676 12628 11732
rect 12572 11340 12628 11396
rect 12908 10722 12964 10724
rect 12908 10670 12910 10722
rect 12910 10670 12962 10722
rect 12962 10670 12964 10722
rect 12908 10668 12964 10670
rect 12460 10108 12516 10164
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 12684 9714 12740 9716
rect 12684 9662 12686 9714
rect 12686 9662 12738 9714
rect 12738 9662 12740 9714
rect 12684 9660 12740 9662
rect 12348 9548 12404 9604
rect 12572 9042 12628 9044
rect 12572 8990 12574 9042
rect 12574 8990 12626 9042
rect 12626 8990 12628 9042
rect 12572 8988 12628 8990
rect 12348 8652 12404 8708
rect 12236 8258 12292 8260
rect 12236 8206 12238 8258
rect 12238 8206 12290 8258
rect 12290 8206 12292 8258
rect 12236 8204 12292 8206
rect 12124 6076 12180 6132
rect 12796 9100 12852 9156
rect 13244 14140 13300 14196
rect 14588 23884 14644 23940
rect 16268 26908 16324 26964
rect 14924 26572 14980 26628
rect 15036 26066 15092 26068
rect 15036 26014 15038 26066
rect 15038 26014 15090 26066
rect 15090 26014 15092 26066
rect 15036 26012 15092 26014
rect 15372 25394 15428 25396
rect 15372 25342 15374 25394
rect 15374 25342 15426 25394
rect 15426 25342 15428 25394
rect 15372 25340 15428 25342
rect 14924 24668 14980 24724
rect 15260 24556 15316 24612
rect 18284 30098 18340 30100
rect 18284 30046 18286 30098
rect 18286 30046 18338 30098
rect 18338 30046 18340 30098
rect 18284 30044 18340 30046
rect 18732 30098 18788 30100
rect 18732 30046 18734 30098
rect 18734 30046 18786 30098
rect 18786 30046 18788 30098
rect 18732 30044 18788 30046
rect 18956 30098 19012 30100
rect 18956 30046 18958 30098
rect 18958 30046 19010 30098
rect 19010 30046 19012 30098
rect 18956 30044 19012 30046
rect 19068 29932 19124 29988
rect 18396 29148 18452 29204
rect 18956 29036 19012 29092
rect 18508 28530 18564 28532
rect 18508 28478 18510 28530
rect 18510 28478 18562 28530
rect 18562 28478 18564 28530
rect 18508 28476 18564 28478
rect 17948 27970 18004 27972
rect 17948 27918 17950 27970
rect 17950 27918 18002 27970
rect 18002 27918 18004 27970
rect 17948 27916 18004 27918
rect 16380 26460 16436 26516
rect 16268 25676 16324 25732
rect 17836 25506 17892 25508
rect 17836 25454 17838 25506
rect 17838 25454 17890 25506
rect 17890 25454 17892 25506
rect 17836 25452 17892 25454
rect 18844 27858 18900 27860
rect 18844 27806 18846 27858
rect 18846 27806 18898 27858
rect 18898 27806 18900 27858
rect 18844 27804 18900 27806
rect 18732 27634 18788 27636
rect 18732 27582 18734 27634
rect 18734 27582 18786 27634
rect 18786 27582 18788 27634
rect 18732 27580 18788 27582
rect 19628 30098 19684 30100
rect 19628 30046 19630 30098
rect 19630 30046 19682 30098
rect 19682 30046 19684 30098
rect 19628 30044 19684 30046
rect 20412 30044 20468 30100
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19180 29148 19236 29204
rect 19068 28924 19124 28980
rect 18732 27132 18788 27188
rect 19068 28476 19124 28532
rect 18396 27074 18452 27076
rect 18396 27022 18398 27074
rect 18398 27022 18450 27074
rect 18450 27022 18452 27074
rect 18396 27020 18452 27022
rect 21756 30828 21812 30884
rect 22316 30882 22372 30884
rect 22316 30830 22318 30882
rect 22318 30830 22370 30882
rect 22370 30830 22372 30882
rect 22316 30828 22372 30830
rect 23436 31218 23492 31220
rect 23436 31166 23438 31218
rect 23438 31166 23490 31218
rect 23490 31166 23492 31218
rect 23436 31164 23492 31166
rect 24780 31388 24836 31444
rect 24444 31218 24500 31220
rect 24444 31166 24446 31218
rect 24446 31166 24498 31218
rect 24498 31166 24500 31218
rect 24444 31164 24500 31166
rect 25340 35698 25396 35700
rect 25340 35646 25342 35698
rect 25342 35646 25394 35698
rect 25394 35646 25396 35698
rect 25340 35644 25396 35646
rect 25564 35308 25620 35364
rect 25452 34690 25508 34692
rect 25452 34638 25454 34690
rect 25454 34638 25506 34690
rect 25506 34638 25508 34690
rect 25452 34636 25508 34638
rect 25452 34076 25508 34132
rect 26012 37996 26068 38052
rect 27020 42588 27076 42644
rect 27132 42364 27188 42420
rect 27468 42812 27524 42868
rect 28028 44940 28084 44996
rect 28140 44882 28196 44884
rect 28140 44830 28142 44882
rect 28142 44830 28194 44882
rect 28194 44830 28196 44882
rect 28140 44828 28196 44830
rect 28252 44322 28308 44324
rect 28252 44270 28254 44322
rect 28254 44270 28306 44322
rect 28306 44270 28308 44322
rect 28252 44268 28308 44270
rect 28140 43260 28196 43316
rect 28140 42866 28196 42868
rect 28140 42814 28142 42866
rect 28142 42814 28194 42866
rect 28194 42814 28196 42866
rect 28140 42812 28196 42814
rect 27468 42530 27524 42532
rect 27468 42478 27470 42530
rect 27470 42478 27522 42530
rect 27522 42478 27524 42530
rect 27468 42476 27524 42478
rect 28140 42588 28196 42644
rect 27356 42140 27412 42196
rect 27468 42252 27524 42308
rect 27020 41244 27076 41300
rect 27916 41916 27972 41972
rect 28028 41692 28084 41748
rect 28140 41356 28196 41412
rect 27580 41244 27636 41300
rect 28028 41186 28084 41188
rect 28028 41134 28030 41186
rect 28030 41134 28082 41186
rect 28082 41134 28084 41186
rect 28028 41132 28084 41134
rect 26572 38780 26628 38836
rect 25900 37938 25956 37940
rect 25900 37886 25902 37938
rect 25902 37886 25954 37938
rect 25954 37886 25956 37938
rect 25900 37884 25956 37886
rect 26012 36482 26068 36484
rect 26012 36430 26014 36482
rect 26014 36430 26066 36482
rect 26066 36430 26068 36482
rect 26012 36428 26068 36430
rect 26348 37660 26404 37716
rect 27356 39900 27412 39956
rect 26684 38892 26740 38948
rect 26908 38444 26964 38500
rect 26684 37660 26740 37716
rect 26796 37324 26852 37380
rect 26908 37212 26964 37268
rect 26572 36540 26628 36596
rect 26796 36204 26852 36260
rect 26572 35868 26628 35924
rect 26236 35196 26292 35252
rect 25788 34914 25844 34916
rect 25788 34862 25790 34914
rect 25790 34862 25842 34914
rect 25842 34862 25844 34914
rect 25788 34860 25844 34862
rect 25900 34524 25956 34580
rect 25676 33740 25732 33796
rect 25788 34412 25844 34468
rect 25676 33570 25732 33572
rect 25676 33518 25678 33570
rect 25678 33518 25730 33570
rect 25730 33518 25732 33570
rect 25676 33516 25732 33518
rect 25340 33458 25396 33460
rect 25340 33406 25342 33458
rect 25342 33406 25394 33458
rect 25394 33406 25396 33458
rect 25340 33404 25396 33406
rect 25228 32844 25284 32900
rect 25452 32732 25508 32788
rect 26012 34188 26068 34244
rect 26124 33964 26180 34020
rect 26348 34076 26404 34132
rect 26684 35308 26740 35364
rect 26684 34914 26740 34916
rect 26684 34862 26686 34914
rect 26686 34862 26738 34914
rect 26738 34862 26740 34914
rect 26684 34860 26740 34862
rect 26684 34412 26740 34468
rect 26684 33852 26740 33908
rect 27916 40402 27972 40404
rect 27916 40350 27918 40402
rect 27918 40350 27970 40402
rect 27970 40350 27972 40402
rect 27916 40348 27972 40350
rect 28140 38834 28196 38836
rect 28140 38782 28142 38834
rect 28142 38782 28194 38834
rect 28194 38782 28196 38834
rect 28140 38780 28196 38782
rect 28700 46620 28756 46676
rect 28588 45106 28644 45108
rect 28588 45054 28590 45106
rect 28590 45054 28642 45106
rect 28642 45054 28644 45106
rect 28588 45052 28644 45054
rect 28588 44716 28644 44772
rect 28588 44380 28644 44436
rect 27804 38444 27860 38500
rect 28588 42530 28644 42532
rect 28588 42478 28590 42530
rect 28590 42478 28642 42530
rect 28642 42478 28644 42530
rect 28588 42476 28644 42478
rect 28476 40460 28532 40516
rect 28700 41804 28756 41860
rect 28700 41244 28756 41300
rect 28588 39900 28644 39956
rect 28476 39730 28532 39732
rect 28476 39678 28478 39730
rect 28478 39678 28530 39730
rect 28530 39678 28532 39730
rect 28476 39676 28532 39678
rect 27916 37884 27972 37940
rect 27468 37324 27524 37380
rect 27356 36876 27412 36932
rect 27020 35868 27076 35924
rect 27020 34636 27076 34692
rect 27356 35644 27412 35700
rect 28252 37548 28308 37604
rect 27916 36482 27972 36484
rect 27916 36430 27918 36482
rect 27918 36430 27970 36482
rect 27970 36430 27972 36482
rect 27916 36428 27972 36430
rect 27580 36204 27636 36260
rect 27468 35084 27524 35140
rect 27132 33628 27188 33684
rect 26908 33068 26964 33124
rect 26572 32844 26628 32900
rect 27580 33180 27636 33236
rect 24892 31164 24948 31220
rect 25116 31388 25172 31444
rect 22764 30882 22820 30884
rect 22764 30830 22766 30882
rect 22766 30830 22818 30882
rect 22818 30830 22820 30882
rect 22764 30828 22820 30830
rect 24668 30882 24724 30884
rect 24668 30830 24670 30882
rect 24670 30830 24722 30882
rect 24722 30830 24724 30882
rect 24668 30828 24724 30830
rect 24332 30268 24388 30324
rect 22988 30098 23044 30100
rect 22988 30046 22990 30098
rect 22990 30046 23042 30098
rect 23042 30046 23044 30098
rect 22988 30044 23044 30046
rect 23660 30044 23716 30100
rect 20972 29932 21028 29988
rect 20636 29372 20692 29428
rect 22092 29426 22148 29428
rect 22092 29374 22094 29426
rect 22094 29374 22146 29426
rect 22146 29374 22148 29426
rect 22092 29372 22148 29374
rect 24556 30156 24612 30212
rect 22540 29036 22596 29092
rect 23548 29148 23604 29204
rect 23212 28700 23268 28756
rect 25452 31666 25508 31668
rect 25452 31614 25454 31666
rect 25454 31614 25506 31666
rect 25506 31614 25508 31666
rect 25452 31612 25508 31614
rect 25340 30882 25396 30884
rect 25340 30830 25342 30882
rect 25342 30830 25394 30882
rect 25394 30830 25396 30882
rect 25340 30828 25396 30830
rect 28924 48242 28980 48244
rect 28924 48190 28926 48242
rect 28926 48190 28978 48242
rect 28978 48190 28980 48242
rect 28924 48188 28980 48190
rect 29036 46562 29092 46564
rect 29036 46510 29038 46562
rect 29038 46510 29090 46562
rect 29090 46510 29092 46562
rect 29036 46508 29092 46510
rect 29260 49308 29316 49364
rect 29932 49196 29988 49252
rect 30044 49026 30100 49028
rect 30044 48974 30046 49026
rect 30046 48974 30098 49026
rect 30098 48974 30100 49026
rect 30044 48972 30100 48974
rect 29932 48188 29988 48244
rect 29260 47458 29316 47460
rect 29260 47406 29262 47458
rect 29262 47406 29314 47458
rect 29314 47406 29316 47458
rect 29260 47404 29316 47406
rect 29596 47404 29652 47460
rect 29260 45778 29316 45780
rect 29260 45726 29262 45778
rect 29262 45726 29314 45778
rect 29314 45726 29316 45778
rect 29260 45724 29316 45726
rect 29148 41468 29204 41524
rect 29484 44380 29540 44436
rect 29708 46060 29764 46116
rect 29932 47570 29988 47572
rect 29932 47518 29934 47570
rect 29934 47518 29986 47570
rect 29986 47518 29988 47570
rect 29932 47516 29988 47518
rect 30716 49810 30772 49812
rect 30716 49758 30718 49810
rect 30718 49758 30770 49810
rect 30770 49758 30772 49810
rect 30716 49756 30772 49758
rect 30380 49084 30436 49140
rect 30604 48972 30660 49028
rect 30828 48748 30884 48804
rect 30268 48636 30324 48692
rect 30156 47682 30212 47684
rect 30156 47630 30158 47682
rect 30158 47630 30210 47682
rect 30210 47630 30212 47682
rect 30156 47628 30212 47630
rect 31164 51436 31220 51492
rect 31164 51266 31220 51268
rect 31164 51214 31166 51266
rect 31166 51214 31218 51266
rect 31218 51214 31220 51266
rect 31164 51212 31220 51214
rect 31388 51100 31444 51156
rect 31052 50316 31108 50372
rect 30604 48524 30660 48580
rect 30828 48242 30884 48244
rect 30828 48190 30830 48242
rect 30830 48190 30882 48242
rect 30882 48190 30884 48242
rect 30828 48188 30884 48190
rect 31052 49420 31108 49476
rect 30828 47292 30884 47348
rect 30828 46674 30884 46676
rect 30828 46622 30830 46674
rect 30830 46622 30882 46674
rect 30882 46622 30884 46674
rect 30828 46620 30884 46622
rect 30492 46562 30548 46564
rect 30492 46510 30494 46562
rect 30494 46510 30546 46562
rect 30546 46510 30548 46562
rect 30492 46508 30548 46510
rect 29932 46060 29988 46116
rect 30156 45836 30212 45892
rect 29708 45666 29764 45668
rect 29708 45614 29710 45666
rect 29710 45614 29762 45666
rect 29762 45614 29764 45666
rect 29708 45612 29764 45614
rect 30044 45778 30100 45780
rect 30044 45726 30046 45778
rect 30046 45726 30098 45778
rect 30098 45726 30100 45778
rect 30044 45724 30100 45726
rect 29708 44716 29764 44772
rect 29708 44156 29764 44212
rect 30604 45666 30660 45668
rect 30604 45614 30606 45666
rect 30606 45614 30658 45666
rect 30658 45614 30660 45666
rect 30604 45612 30660 45614
rect 29932 44268 29988 44324
rect 31500 50316 31556 50372
rect 31276 49308 31332 49364
rect 31388 48802 31444 48804
rect 31388 48750 31390 48802
rect 31390 48750 31442 48802
rect 31442 48750 31444 48802
rect 31388 48748 31444 48750
rect 31164 47404 31220 47460
rect 33516 55970 33572 55972
rect 33516 55918 33518 55970
rect 33518 55918 33570 55970
rect 33570 55918 33572 55970
rect 33516 55916 33572 55918
rect 31948 54572 32004 54628
rect 31948 53676 32004 53732
rect 32284 52834 32340 52836
rect 32284 52782 32286 52834
rect 32286 52782 32338 52834
rect 32338 52782 32340 52834
rect 32284 52780 32340 52782
rect 31724 52668 31780 52724
rect 31836 50482 31892 50484
rect 31836 50430 31838 50482
rect 31838 50430 31890 50482
rect 31890 50430 31892 50482
rect 31836 50428 31892 50430
rect 31612 49420 31668 49476
rect 31612 49084 31668 49140
rect 32172 48466 32228 48468
rect 32172 48414 32174 48466
rect 32174 48414 32226 48466
rect 32226 48414 32228 48466
rect 32172 48412 32228 48414
rect 32060 48242 32116 48244
rect 32060 48190 32062 48242
rect 32062 48190 32114 48242
rect 32114 48190 32116 48242
rect 32060 48188 32116 48190
rect 31164 47234 31220 47236
rect 31164 47182 31166 47234
rect 31166 47182 31218 47234
rect 31218 47182 31220 47234
rect 31164 47180 31220 47182
rect 31276 46956 31332 47012
rect 31500 47292 31556 47348
rect 31164 46508 31220 46564
rect 31164 45724 31220 45780
rect 29260 41692 29316 41748
rect 29148 40796 29204 40852
rect 29372 40572 29428 40628
rect 29260 40124 29316 40180
rect 29596 40124 29652 40180
rect 29372 39564 29428 39620
rect 29372 39340 29428 39396
rect 29596 39058 29652 39060
rect 29596 39006 29598 39058
rect 29598 39006 29650 39058
rect 29650 39006 29652 39058
rect 29596 39004 29652 39006
rect 29148 38946 29204 38948
rect 29148 38894 29150 38946
rect 29150 38894 29202 38946
rect 29202 38894 29204 38946
rect 29148 38892 29204 38894
rect 28364 36876 28420 36932
rect 28140 35026 28196 35028
rect 28140 34974 28142 35026
rect 28142 34974 28194 35026
rect 28194 34974 28196 35026
rect 28140 34972 28196 34974
rect 28140 33458 28196 33460
rect 28140 33406 28142 33458
rect 28142 33406 28194 33458
rect 28194 33406 28196 33458
rect 28140 33404 28196 33406
rect 29820 40572 29876 40628
rect 29260 37938 29316 37940
rect 29260 37886 29262 37938
rect 29262 37886 29314 37938
rect 29314 37886 29316 37938
rect 29260 37884 29316 37886
rect 29372 37660 29428 37716
rect 29260 36594 29316 36596
rect 29260 36542 29262 36594
rect 29262 36542 29314 36594
rect 29314 36542 29316 36594
rect 29260 36540 29316 36542
rect 29036 35922 29092 35924
rect 29036 35870 29038 35922
rect 29038 35870 29090 35922
rect 29090 35870 29092 35922
rect 29036 35868 29092 35870
rect 28924 35698 28980 35700
rect 28924 35646 28926 35698
rect 28926 35646 28978 35698
rect 28978 35646 28980 35698
rect 28924 35644 28980 35646
rect 28364 35308 28420 35364
rect 28476 35084 28532 35140
rect 29260 35308 29316 35364
rect 29260 34972 29316 35028
rect 29148 34860 29204 34916
rect 28476 34802 28532 34804
rect 28476 34750 28478 34802
rect 28478 34750 28530 34802
rect 28530 34750 28532 34802
rect 28476 34748 28532 34750
rect 29036 34130 29092 34132
rect 29036 34078 29038 34130
rect 29038 34078 29090 34130
rect 29090 34078 29092 34130
rect 29036 34076 29092 34078
rect 28700 33852 28756 33908
rect 28364 33404 28420 33460
rect 28476 33180 28532 33236
rect 28140 32956 28196 33012
rect 29484 34914 29540 34916
rect 29484 34862 29486 34914
rect 29486 34862 29538 34914
rect 29538 34862 29540 34914
rect 29484 34860 29540 34862
rect 30492 44492 30548 44548
rect 30604 44268 30660 44324
rect 30940 44940 30996 44996
rect 30492 43372 30548 43428
rect 30380 42642 30436 42644
rect 30380 42590 30382 42642
rect 30382 42590 30434 42642
rect 30434 42590 30436 42642
rect 30380 42588 30436 42590
rect 30268 41970 30324 41972
rect 30268 41918 30270 41970
rect 30270 41918 30322 41970
rect 30322 41918 30324 41970
rect 30268 41916 30324 41918
rect 30604 42812 30660 42868
rect 30940 44268 30996 44324
rect 31500 46060 31556 46116
rect 31388 44882 31444 44884
rect 31388 44830 31390 44882
rect 31390 44830 31442 44882
rect 31442 44830 31444 44882
rect 31388 44828 31444 44830
rect 31612 45890 31668 45892
rect 31612 45838 31614 45890
rect 31614 45838 31666 45890
rect 31666 45838 31668 45890
rect 31612 45836 31668 45838
rect 31836 45778 31892 45780
rect 31836 45726 31838 45778
rect 31838 45726 31890 45778
rect 31890 45726 31892 45778
rect 31836 45724 31892 45726
rect 31836 45388 31892 45444
rect 32620 47180 32676 47236
rect 32508 45948 32564 46004
rect 33068 55298 33124 55300
rect 33068 55246 33070 55298
rect 33070 55246 33122 55298
rect 33122 55246 33124 55298
rect 33068 55244 33124 55246
rect 33180 54626 33236 54628
rect 33180 54574 33182 54626
rect 33182 54574 33234 54626
rect 33234 54574 33236 54626
rect 33180 54572 33236 54574
rect 32956 52892 33012 52948
rect 33292 53564 33348 53620
rect 34076 55298 34132 55300
rect 34076 55246 34078 55298
rect 34078 55246 34130 55298
rect 34130 55246 34132 55298
rect 34076 55244 34132 55246
rect 33852 55132 33908 55188
rect 34860 55916 34916 55972
rect 33852 54684 33908 54740
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 48972 56306 49028 56308
rect 48972 56254 48974 56306
rect 48974 56254 49026 56306
rect 49026 56254 49028 56306
rect 48972 56252 49028 56254
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 49196 56252 49252 56308
rect 48412 55356 48468 55412
rect 49532 56028 49588 56084
rect 34076 54348 34132 54404
rect 33852 54236 33908 54292
rect 34412 53730 34468 53732
rect 34412 53678 34414 53730
rect 34414 53678 34466 53730
rect 34466 53678 34468 53730
rect 34412 53676 34468 53678
rect 33180 51100 33236 51156
rect 32956 50482 33012 50484
rect 32956 50430 32958 50482
rect 32958 50430 33010 50482
rect 33010 50430 33012 50482
rect 32956 50428 33012 50430
rect 33292 50594 33348 50596
rect 33292 50542 33294 50594
rect 33294 50542 33346 50594
rect 33346 50542 33348 50594
rect 33292 50540 33348 50542
rect 33292 48972 33348 49028
rect 33068 48748 33124 48804
rect 31948 44940 32004 44996
rect 32284 44268 32340 44324
rect 30716 42700 30772 42756
rect 30268 39900 30324 39956
rect 30940 42028 30996 42084
rect 31388 42642 31444 42644
rect 31388 42590 31390 42642
rect 31390 42590 31442 42642
rect 31442 42590 31444 42642
rect 31388 42588 31444 42590
rect 31612 42530 31668 42532
rect 31612 42478 31614 42530
rect 31614 42478 31666 42530
rect 31666 42478 31668 42530
rect 31612 42476 31668 42478
rect 30940 40796 30996 40852
rect 31052 40124 31108 40180
rect 30492 40012 30548 40068
rect 30268 39564 30324 39620
rect 30380 39340 30436 39396
rect 29820 36988 29876 37044
rect 30268 37154 30324 37156
rect 30268 37102 30270 37154
rect 30270 37102 30322 37154
rect 30322 37102 30324 37154
rect 30268 37100 30324 37102
rect 30604 38892 30660 38948
rect 31612 40908 31668 40964
rect 31500 40572 31556 40628
rect 32284 43538 32340 43540
rect 32284 43486 32286 43538
rect 32286 43486 32338 43538
rect 32338 43486 32340 43538
rect 32284 43484 32340 43486
rect 31948 43426 32004 43428
rect 31948 43374 31950 43426
rect 31950 43374 32002 43426
rect 32002 43374 32004 43426
rect 31948 43372 32004 43374
rect 32620 43372 32676 43428
rect 32172 42364 32228 42420
rect 32172 41356 32228 41412
rect 32396 41298 32452 41300
rect 32396 41246 32398 41298
rect 32398 41246 32450 41298
rect 32450 41246 32452 41298
rect 32396 41244 32452 41246
rect 32508 41804 32564 41860
rect 32172 40572 32228 40628
rect 30828 39788 30884 39844
rect 31388 39618 31444 39620
rect 31388 39566 31390 39618
rect 31390 39566 31442 39618
rect 31442 39566 31444 39618
rect 31388 39564 31444 39566
rect 31164 39452 31220 39508
rect 31388 39228 31444 39284
rect 30940 38892 30996 38948
rect 30828 38780 30884 38836
rect 31612 40124 31668 40180
rect 31612 39900 31668 39956
rect 31612 38834 31668 38836
rect 31612 38782 31614 38834
rect 31614 38782 31666 38834
rect 31666 38782 31668 38834
rect 31612 38780 31668 38782
rect 30716 37660 30772 37716
rect 31500 38220 31556 38276
rect 31836 40178 31892 40180
rect 31836 40126 31838 40178
rect 31838 40126 31890 40178
rect 31890 40126 31892 40178
rect 31836 40124 31892 40126
rect 31612 38108 31668 38164
rect 31948 37938 32004 37940
rect 31948 37886 31950 37938
rect 31950 37886 32002 37938
rect 32002 37886 32004 37938
rect 31948 37884 32004 37886
rect 30716 37154 30772 37156
rect 30716 37102 30718 37154
rect 30718 37102 30770 37154
rect 30770 37102 30772 37154
rect 30716 37100 30772 37102
rect 30156 36428 30212 36484
rect 30268 35980 30324 36036
rect 29820 35532 29876 35588
rect 29820 33964 29876 34020
rect 29708 33068 29764 33124
rect 30044 35420 30100 35476
rect 30604 36204 30660 36260
rect 30604 35586 30660 35588
rect 30604 35534 30606 35586
rect 30606 35534 30658 35586
rect 30658 35534 30660 35586
rect 30604 35532 30660 35534
rect 30380 34748 30436 34804
rect 30940 36428 30996 36484
rect 31052 36876 31108 36932
rect 30940 36204 30996 36260
rect 30940 35980 30996 36036
rect 31612 37100 31668 37156
rect 31500 36876 31556 36932
rect 32284 38162 32340 38164
rect 32284 38110 32286 38162
rect 32286 38110 32338 38162
rect 32338 38110 32340 38162
rect 32284 38108 32340 38110
rect 32172 36764 32228 36820
rect 32396 37100 32452 37156
rect 32620 38050 32676 38052
rect 32620 37998 32622 38050
rect 32622 37998 32674 38050
rect 32674 37998 32676 38050
rect 32620 37996 32676 37998
rect 32844 45890 32900 45892
rect 32844 45838 32846 45890
rect 32846 45838 32898 45890
rect 32898 45838 32900 45890
rect 32844 45836 32900 45838
rect 32844 45388 32900 45444
rect 34076 52780 34132 52836
rect 34300 52892 34356 52948
rect 36988 55298 37044 55300
rect 36988 55246 36990 55298
rect 36990 55246 37042 55298
rect 37042 55246 37044 55298
rect 36988 55244 37044 55246
rect 35420 54348 35476 54404
rect 35196 54236 35252 54292
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35084 53564 35140 53620
rect 36092 53676 36148 53732
rect 35868 53564 35924 53620
rect 34748 52946 34804 52948
rect 34748 52894 34750 52946
rect 34750 52894 34802 52946
rect 34802 52894 34804 52946
rect 34748 52892 34804 52894
rect 34972 52892 35028 52948
rect 34636 52834 34692 52836
rect 34636 52782 34638 52834
rect 34638 52782 34690 52834
rect 34690 52782 34692 52834
rect 34636 52780 34692 52782
rect 34860 52332 34916 52388
rect 34076 51266 34132 51268
rect 34076 51214 34078 51266
rect 34078 51214 34130 51266
rect 34130 51214 34132 51266
rect 34076 51212 34132 51214
rect 34748 51154 34804 51156
rect 34748 51102 34750 51154
rect 34750 51102 34802 51154
rect 34802 51102 34804 51154
rect 34748 51100 34804 51102
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35084 52108 35140 52164
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 33964 50594 34020 50596
rect 33964 50542 33966 50594
rect 33966 50542 34018 50594
rect 34018 50542 34020 50594
rect 33964 50540 34020 50542
rect 35420 50034 35476 50036
rect 35420 49982 35422 50034
rect 35422 49982 35474 50034
rect 35474 49982 35476 50034
rect 35420 49980 35476 49982
rect 35644 49756 35700 49812
rect 33852 48188 33908 48244
rect 34076 49026 34132 49028
rect 34076 48974 34078 49026
rect 34078 48974 34130 49026
rect 34130 48974 34132 49026
rect 34076 48972 34132 48974
rect 35420 49644 35476 49700
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34524 49084 34580 49140
rect 34076 48188 34132 48244
rect 33404 47628 33460 47684
rect 33628 47740 33684 47796
rect 33516 45890 33572 45892
rect 33516 45838 33518 45890
rect 33518 45838 33570 45890
rect 33570 45838 33572 45890
rect 33516 45836 33572 45838
rect 33740 45778 33796 45780
rect 33740 45726 33742 45778
rect 33742 45726 33794 45778
rect 33794 45726 33796 45778
rect 33740 45724 33796 45726
rect 34300 47628 34356 47684
rect 35420 48412 35476 48468
rect 35532 48972 35588 49028
rect 36428 53506 36484 53508
rect 36428 53454 36430 53506
rect 36430 53454 36482 53506
rect 36482 53454 36484 53506
rect 36428 53452 36484 53454
rect 36316 52892 36372 52948
rect 37772 54348 37828 54404
rect 37996 53842 38052 53844
rect 37996 53790 37998 53842
rect 37998 53790 38050 53842
rect 38050 53790 38052 53842
rect 37996 53788 38052 53790
rect 37324 53676 37380 53732
rect 37212 53564 37268 53620
rect 38444 54402 38500 54404
rect 38444 54350 38446 54402
rect 38446 54350 38498 54402
rect 38498 54350 38500 54402
rect 38444 54348 38500 54350
rect 38108 53564 38164 53620
rect 36092 51378 36148 51380
rect 36092 51326 36094 51378
rect 36094 51326 36146 51378
rect 36146 51326 36148 51378
rect 36092 51324 36148 51326
rect 37100 52892 37156 52948
rect 41020 55186 41076 55188
rect 41020 55134 41022 55186
rect 41022 55134 41074 55186
rect 41074 55134 41076 55186
rect 41020 55132 41076 55134
rect 42476 55186 42532 55188
rect 42476 55134 42478 55186
rect 42478 55134 42530 55186
rect 42530 55134 42532 55186
rect 42476 55132 42532 55134
rect 39900 54348 39956 54404
rect 39788 53900 39844 53956
rect 41356 53842 41412 53844
rect 41356 53790 41358 53842
rect 41358 53790 41410 53842
rect 41410 53790 41412 53842
rect 41356 53788 41412 53790
rect 39452 53618 39508 53620
rect 39452 53566 39454 53618
rect 39454 53566 39506 53618
rect 39506 53566 39508 53618
rect 39452 53564 39508 53566
rect 42140 55074 42196 55076
rect 42140 55022 42142 55074
rect 42142 55022 42194 55074
rect 42194 55022 42196 55074
rect 42140 55020 42196 55022
rect 42252 54514 42308 54516
rect 42252 54462 42254 54514
rect 42254 54462 42306 54514
rect 42306 54462 42308 54514
rect 42252 54460 42308 54462
rect 38108 52332 38164 52388
rect 38444 52668 38500 52724
rect 42924 55132 42980 55188
rect 42588 54236 42644 54292
rect 42028 53452 42084 53508
rect 37548 51884 37604 51940
rect 36988 51490 37044 51492
rect 36988 51438 36990 51490
rect 36990 51438 37042 51490
rect 37042 51438 37044 51490
rect 36988 51436 37044 51438
rect 37548 50540 37604 50596
rect 37660 51100 37716 51156
rect 36876 50204 36932 50260
rect 36428 49756 36484 49812
rect 35644 48748 35700 48804
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 36540 48748 36596 48804
rect 36540 48242 36596 48244
rect 36540 48190 36542 48242
rect 36542 48190 36594 48242
rect 36594 48190 36596 48242
rect 36540 48188 36596 48190
rect 36316 47628 36372 47684
rect 34300 45948 34356 46004
rect 34636 45948 34692 46004
rect 34412 45106 34468 45108
rect 34412 45054 34414 45106
rect 34414 45054 34466 45106
rect 34466 45054 34468 45106
rect 34412 45052 34468 45054
rect 34524 45724 34580 45780
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 46002 35252 46004
rect 35196 45950 35198 46002
rect 35198 45950 35250 46002
rect 35250 45950 35252 46002
rect 35196 45948 35252 45950
rect 35084 45890 35140 45892
rect 35084 45838 35086 45890
rect 35086 45838 35138 45890
rect 35138 45838 35140 45890
rect 35084 45836 35140 45838
rect 34188 44940 34244 44996
rect 33852 43484 33908 43540
rect 33740 42028 33796 42084
rect 33180 41858 33236 41860
rect 33180 41806 33182 41858
rect 33182 41806 33234 41858
rect 33234 41806 33236 41858
rect 33180 41804 33236 41806
rect 33516 41580 33572 41636
rect 33516 41244 33572 41300
rect 33292 40684 33348 40740
rect 33180 40572 33236 40628
rect 32956 39004 33012 39060
rect 33516 40460 33572 40516
rect 33404 38556 33460 38612
rect 32844 38220 32900 38276
rect 34300 44604 34356 44660
rect 34300 43036 34356 43092
rect 34300 42866 34356 42868
rect 34300 42814 34302 42866
rect 34302 42814 34354 42866
rect 34354 42814 34356 42866
rect 34300 42812 34356 42814
rect 34300 42252 34356 42308
rect 34412 42082 34468 42084
rect 34412 42030 34414 42082
rect 34414 42030 34466 42082
rect 34466 42030 34468 42082
rect 34412 42028 34468 42030
rect 34300 41804 34356 41860
rect 34412 41074 34468 41076
rect 34412 41022 34414 41074
rect 34414 41022 34466 41074
rect 34466 41022 34468 41074
rect 34412 41020 34468 41022
rect 34748 43484 34804 43540
rect 34972 43036 35028 43092
rect 34860 42812 34916 42868
rect 34748 42140 34804 42196
rect 34636 41916 34692 41972
rect 35196 44994 35252 44996
rect 35196 44942 35198 44994
rect 35198 44942 35250 44994
rect 35250 44942 35252 44994
rect 35196 44940 35252 44942
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35308 44322 35364 44324
rect 35308 44270 35310 44322
rect 35310 44270 35362 44322
rect 35362 44270 35364 44322
rect 35308 44268 35364 44270
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34300 40514 34356 40516
rect 34300 40462 34302 40514
rect 34302 40462 34354 40514
rect 34354 40462 34356 40514
rect 34300 40460 34356 40462
rect 34076 40348 34132 40404
rect 34188 39842 34244 39844
rect 34188 39790 34190 39842
rect 34190 39790 34242 39842
rect 34242 39790 34244 39842
rect 34188 39788 34244 39790
rect 34860 40236 34916 40292
rect 35308 42364 35364 42420
rect 35308 41970 35364 41972
rect 35308 41918 35310 41970
rect 35310 41918 35362 41970
rect 35362 41918 35364 41970
rect 35308 41916 35364 41918
rect 36540 47458 36596 47460
rect 36540 47406 36542 47458
rect 36542 47406 36594 47458
rect 36594 47406 36596 47458
rect 36540 47404 36596 47406
rect 35868 46114 35924 46116
rect 35868 46062 35870 46114
rect 35870 46062 35922 46114
rect 35922 46062 35924 46114
rect 35868 46060 35924 46062
rect 35644 42642 35700 42644
rect 35644 42590 35646 42642
rect 35646 42590 35698 42642
rect 35698 42590 35700 42642
rect 35644 42588 35700 42590
rect 36316 47234 36372 47236
rect 36316 47182 36318 47234
rect 36318 47182 36370 47234
rect 36370 47182 36372 47234
rect 36316 47180 36372 47182
rect 37212 47458 37268 47460
rect 37212 47406 37214 47458
rect 37214 47406 37266 47458
rect 37266 47406 37268 47458
rect 37212 47404 37268 47406
rect 37100 47180 37156 47236
rect 36988 44322 37044 44324
rect 36988 44270 36990 44322
rect 36990 44270 37042 44322
rect 37042 44270 37044 44322
rect 36988 44268 37044 44270
rect 37884 51154 37940 51156
rect 37884 51102 37886 51154
rect 37886 51102 37938 51154
rect 37938 51102 37940 51154
rect 37884 51100 37940 51102
rect 38780 51996 38836 52052
rect 38556 51324 38612 51380
rect 38332 50652 38388 50708
rect 38780 51100 38836 51156
rect 39452 51938 39508 51940
rect 39452 51886 39454 51938
rect 39454 51886 39506 51938
rect 39506 51886 39508 51938
rect 39452 51884 39508 51886
rect 39004 50652 39060 50708
rect 39116 51378 39172 51380
rect 39116 51326 39118 51378
rect 39118 51326 39170 51378
rect 39170 51326 39172 51378
rect 39116 51324 39172 51326
rect 39004 50482 39060 50484
rect 39004 50430 39006 50482
rect 39006 50430 39058 50482
rect 39058 50430 39060 50482
rect 39004 50428 39060 50430
rect 40012 51324 40068 51380
rect 40796 51938 40852 51940
rect 40796 51886 40798 51938
rect 40798 51886 40850 51938
rect 40850 51886 40852 51938
rect 40796 51884 40852 51886
rect 41020 51660 41076 51716
rect 39228 51100 39284 51156
rect 39788 50652 39844 50708
rect 39340 50594 39396 50596
rect 39340 50542 39342 50594
rect 39342 50542 39394 50594
rect 39394 50542 39396 50594
rect 39340 50540 39396 50542
rect 38108 50034 38164 50036
rect 38108 49982 38110 50034
rect 38110 49982 38162 50034
rect 38162 49982 38164 50034
rect 38108 49980 38164 49982
rect 37660 49868 37716 49924
rect 37436 49644 37492 49700
rect 37996 49698 38052 49700
rect 37996 49646 37998 49698
rect 37998 49646 38050 49698
rect 38050 49646 38052 49698
rect 37996 49644 38052 49646
rect 37884 48972 37940 49028
rect 38444 48972 38500 49028
rect 39004 49138 39060 49140
rect 39004 49086 39006 49138
rect 39006 49086 39058 49138
rect 39058 49086 39060 49138
rect 39004 49084 39060 49086
rect 39004 48748 39060 48804
rect 37436 47628 37492 47684
rect 37660 47516 37716 47572
rect 37324 44546 37380 44548
rect 37324 44494 37326 44546
rect 37326 44494 37378 44546
rect 37378 44494 37380 44546
rect 37324 44492 37380 44494
rect 36316 43484 36372 43540
rect 35868 42812 35924 42868
rect 35756 42364 35812 42420
rect 35980 42140 36036 42196
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35084 41074 35140 41076
rect 35084 41022 35086 41074
rect 35086 41022 35138 41074
rect 35138 41022 35140 41074
rect 35084 41020 35140 41022
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35084 39788 35140 39844
rect 36316 40290 36372 40292
rect 36316 40238 36318 40290
rect 36318 40238 36370 40290
rect 36370 40238 36372 40290
rect 36316 40236 36372 40238
rect 36428 39506 36484 39508
rect 36428 39454 36430 39506
rect 36430 39454 36482 39506
rect 36482 39454 36484 39506
rect 36428 39452 36484 39454
rect 32732 37772 32788 37828
rect 33180 37212 33236 37268
rect 33964 37884 34020 37940
rect 33740 36988 33796 37044
rect 33516 36652 33572 36708
rect 32508 36316 32564 36372
rect 32060 35980 32116 36036
rect 31724 35810 31780 35812
rect 31724 35758 31726 35810
rect 31726 35758 31778 35810
rect 31778 35758 31780 35810
rect 31724 35756 31780 35758
rect 31388 35644 31444 35700
rect 31276 35196 31332 35252
rect 33068 36482 33124 36484
rect 33068 36430 33070 36482
rect 33070 36430 33122 36482
rect 33122 36430 33124 36482
rect 33068 36428 33124 36430
rect 33852 35868 33908 35924
rect 33628 35420 33684 35476
rect 32732 35196 32788 35252
rect 31948 34972 32004 35028
rect 31164 34860 31220 34916
rect 30716 34524 30772 34580
rect 31164 34524 31220 34580
rect 30716 33964 30772 34020
rect 30940 33346 30996 33348
rect 30940 33294 30942 33346
rect 30942 33294 30994 33346
rect 30994 33294 30996 33346
rect 30940 33292 30996 33294
rect 30380 32786 30436 32788
rect 30380 32734 30382 32786
rect 30382 32734 30434 32786
rect 30434 32734 30436 32786
rect 30380 32732 30436 32734
rect 28028 31724 28084 31780
rect 25116 30268 25172 30324
rect 25004 30044 25060 30100
rect 24444 29986 24500 29988
rect 24444 29934 24446 29986
rect 24446 29934 24498 29986
rect 24498 29934 24500 29986
rect 24444 29932 24500 29934
rect 25452 30156 25508 30212
rect 25116 29986 25172 29988
rect 25116 29934 25118 29986
rect 25118 29934 25170 29986
rect 25170 29934 25172 29986
rect 25116 29932 25172 29934
rect 24332 29148 24388 29204
rect 24668 29036 24724 29092
rect 23772 28700 23828 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 28028 19684 28084
rect 25004 28642 25060 28644
rect 25004 28590 25006 28642
rect 25006 28590 25058 28642
rect 25058 28590 25060 28642
rect 25004 28588 25060 28590
rect 25788 30098 25844 30100
rect 25788 30046 25790 30098
rect 25790 30046 25842 30098
rect 25842 30046 25844 30098
rect 25788 30044 25844 30046
rect 25900 28700 25956 28756
rect 25564 28588 25620 28644
rect 24668 28082 24724 28084
rect 24668 28030 24670 28082
rect 24670 28030 24722 28082
rect 24722 28030 24724 28082
rect 24668 28028 24724 28030
rect 25676 28364 25732 28420
rect 19404 27916 19460 27972
rect 21756 27692 21812 27748
rect 18172 25452 18228 25508
rect 16044 25394 16100 25396
rect 16044 25342 16046 25394
rect 16046 25342 16098 25394
rect 16098 25342 16100 25394
rect 16044 25340 16100 25342
rect 16604 25228 16660 25284
rect 15484 24892 15540 24948
rect 16268 23436 16324 23492
rect 14588 22370 14644 22372
rect 14588 22318 14590 22370
rect 14590 22318 14642 22370
rect 14642 22318 14644 22370
rect 14588 22316 14644 22318
rect 14476 21420 14532 21476
rect 14700 21474 14756 21476
rect 14700 21422 14702 21474
rect 14702 21422 14754 21474
rect 14754 21422 14756 21474
rect 14700 21420 14756 21422
rect 14812 20300 14868 20356
rect 14588 19852 14644 19908
rect 14476 19740 14532 19796
rect 14364 17500 14420 17556
rect 13916 17388 13972 17444
rect 13804 16940 13860 16996
rect 16268 23154 16324 23156
rect 16268 23102 16270 23154
rect 16270 23102 16322 23154
rect 16322 23102 16324 23154
rect 16268 23100 16324 23102
rect 15372 22428 15428 22484
rect 15148 22258 15204 22260
rect 15148 22206 15150 22258
rect 15150 22206 15202 22258
rect 15202 22206 15204 22258
rect 15148 22204 15204 22206
rect 15820 22204 15876 22260
rect 15484 21644 15540 21700
rect 15148 21586 15204 21588
rect 15148 21534 15150 21586
rect 15150 21534 15202 21586
rect 15202 21534 15204 21586
rect 15148 21532 15204 21534
rect 15484 20188 15540 20244
rect 15148 19404 15204 19460
rect 14812 18450 14868 18452
rect 14812 18398 14814 18450
rect 14814 18398 14866 18450
rect 14866 18398 14868 18450
rect 14812 18396 14868 18398
rect 14588 17948 14644 18004
rect 14700 17724 14756 17780
rect 14588 16828 14644 16884
rect 13804 16770 13860 16772
rect 13804 16718 13806 16770
rect 13806 16718 13858 16770
rect 13858 16718 13860 16770
rect 13804 16716 13860 16718
rect 14140 16716 14196 16772
rect 14140 16492 14196 16548
rect 13692 15596 13748 15652
rect 15036 17052 15092 17108
rect 13468 14588 13524 14644
rect 13804 15036 13860 15092
rect 13692 14364 13748 14420
rect 13580 12460 13636 12516
rect 13804 14252 13860 14308
rect 13692 11564 13748 11620
rect 13244 10556 13300 10612
rect 13804 10892 13860 10948
rect 13132 9548 13188 9604
rect 12908 8428 12964 8484
rect 12796 8092 12852 8148
rect 13356 10108 13412 10164
rect 13356 8930 13412 8932
rect 13356 8878 13358 8930
rect 13358 8878 13410 8930
rect 13410 8878 13412 8930
rect 13356 8876 13412 8878
rect 13692 9884 13748 9940
rect 14812 16044 14868 16100
rect 14028 13692 14084 13748
rect 14028 11788 14084 11844
rect 14028 11004 14084 11060
rect 14028 10668 14084 10724
rect 13916 10332 13972 10388
rect 13580 9660 13636 9716
rect 13692 9324 13748 9380
rect 13692 8988 13748 9044
rect 13580 8428 13636 8484
rect 13580 8204 13636 8260
rect 13804 7980 13860 8036
rect 13244 7644 13300 7700
rect 12684 6524 12740 6580
rect 12572 6076 12628 6132
rect 12124 5852 12180 5908
rect 11564 5234 11620 5236
rect 11564 5182 11566 5234
rect 11566 5182 11618 5234
rect 11618 5182 11620 5234
rect 11564 5180 11620 5182
rect 11788 4956 11844 5012
rect 11564 3612 11620 3668
rect 10780 3276 10836 3332
rect 8988 3164 9044 3220
rect 8316 2828 8372 2884
rect 11900 4450 11956 4452
rect 11900 4398 11902 4450
rect 11902 4398 11954 4450
rect 11954 4398 11956 4450
rect 11900 4396 11956 4398
rect 13020 7420 13076 7476
rect 13132 7532 13188 7588
rect 12908 6860 12964 6916
rect 13244 6748 13300 6804
rect 13356 7756 13412 7812
rect 14812 15596 14868 15652
rect 14588 15484 14644 15540
rect 14476 15036 14532 15092
rect 14476 14252 14532 14308
rect 14588 13916 14644 13972
rect 14700 13746 14756 13748
rect 14700 13694 14702 13746
rect 14702 13694 14754 13746
rect 14754 13694 14756 13746
rect 14700 13692 14756 13694
rect 14252 13020 14308 13076
rect 14476 13020 14532 13076
rect 14364 12962 14420 12964
rect 14364 12910 14366 12962
rect 14366 12910 14418 12962
rect 14418 12910 14420 12962
rect 14364 12908 14420 12910
rect 14252 10220 14308 10276
rect 14588 12684 14644 12740
rect 17388 24722 17444 24724
rect 17388 24670 17390 24722
rect 17390 24670 17442 24722
rect 17442 24670 17444 24722
rect 17388 24668 17444 24670
rect 16492 23938 16548 23940
rect 16492 23886 16494 23938
rect 16494 23886 16546 23938
rect 16546 23886 16548 23938
rect 16492 23884 16548 23886
rect 16492 23548 16548 23604
rect 18732 25506 18788 25508
rect 18732 25454 18734 25506
rect 18734 25454 18786 25506
rect 18786 25454 18788 25506
rect 18732 25452 18788 25454
rect 17836 24892 17892 24948
rect 17612 24332 17668 24388
rect 18060 24332 18116 24388
rect 16716 23212 16772 23268
rect 16044 21980 16100 22036
rect 16380 22370 16436 22372
rect 16380 22318 16382 22370
rect 16382 22318 16434 22370
rect 16434 22318 16436 22370
rect 16380 22316 16436 22318
rect 17164 22428 17220 22484
rect 16716 21868 16772 21924
rect 16492 21756 16548 21812
rect 16044 21532 16100 21588
rect 15596 19404 15652 19460
rect 15708 20188 15764 20244
rect 15260 17612 15316 17668
rect 15148 16044 15204 16100
rect 15708 17948 15764 18004
rect 15036 15932 15092 15988
rect 15036 15372 15092 15428
rect 15484 16828 15540 16884
rect 15372 16156 15428 16212
rect 15372 15596 15428 15652
rect 14924 14476 14980 14532
rect 15820 17666 15876 17668
rect 15820 17614 15822 17666
rect 15822 17614 15874 17666
rect 15874 17614 15876 17666
rect 15820 17612 15876 17614
rect 15820 17276 15876 17332
rect 15596 16492 15652 16548
rect 15596 15484 15652 15540
rect 15820 16098 15876 16100
rect 15820 16046 15822 16098
rect 15822 16046 15874 16098
rect 15874 16046 15876 16098
rect 15820 16044 15876 16046
rect 14924 13468 14980 13524
rect 15372 14642 15428 14644
rect 15372 14590 15374 14642
rect 15374 14590 15426 14642
rect 15426 14590 15428 14642
rect 15372 14588 15428 14590
rect 15372 14028 15428 14084
rect 15260 13468 15316 13524
rect 15596 13916 15652 13972
rect 15484 13468 15540 13524
rect 15036 12962 15092 12964
rect 15036 12910 15038 12962
rect 15038 12910 15090 12962
rect 15090 12910 15092 12962
rect 15036 12908 15092 12910
rect 14140 10108 14196 10164
rect 14364 9996 14420 10052
rect 14588 11676 14644 11732
rect 14588 10332 14644 10388
rect 14700 11228 14756 11284
rect 14924 11676 14980 11732
rect 14812 10892 14868 10948
rect 15596 12236 15652 12292
rect 15036 11004 15092 11060
rect 14924 10556 14980 10612
rect 14924 10220 14980 10276
rect 14812 10108 14868 10164
rect 14476 9772 14532 9828
rect 13916 7532 13972 7588
rect 14588 9660 14644 9716
rect 13468 7474 13524 7476
rect 13468 7422 13470 7474
rect 13470 7422 13522 7474
rect 13522 7422 13524 7474
rect 13468 7420 13524 7422
rect 13692 7250 13748 7252
rect 13692 7198 13694 7250
rect 13694 7198 13746 7250
rect 13746 7198 13748 7250
rect 13692 7196 13748 7198
rect 12908 6412 12964 6468
rect 12684 5292 12740 5348
rect 13356 6524 13412 6580
rect 14140 9154 14196 9156
rect 14140 9102 14142 9154
rect 14142 9102 14194 9154
rect 14194 9102 14196 9154
rect 14140 9100 14196 9102
rect 14476 8316 14532 8372
rect 14700 8370 14756 8372
rect 14700 8318 14702 8370
rect 14702 8318 14754 8370
rect 14754 8318 14756 8370
rect 14700 8316 14756 8318
rect 15260 10332 15316 10388
rect 15372 9996 15428 10052
rect 15372 9772 15428 9828
rect 15484 9660 15540 9716
rect 15260 9436 15316 9492
rect 14924 9042 14980 9044
rect 14924 8990 14926 9042
rect 14926 8990 14978 9042
rect 14978 8990 14980 9042
rect 14924 8988 14980 8990
rect 15484 8764 15540 8820
rect 15372 8540 15428 8596
rect 14140 8092 14196 8148
rect 13244 5180 13300 5236
rect 12236 5122 12292 5124
rect 12236 5070 12238 5122
rect 12238 5070 12290 5122
rect 12290 5070 12292 5122
rect 12236 5068 12292 5070
rect 13468 5346 13524 5348
rect 13468 5294 13470 5346
rect 13470 5294 13522 5346
rect 13522 5294 13524 5346
rect 13468 5292 13524 5294
rect 14028 6690 14084 6692
rect 14028 6638 14030 6690
rect 14030 6638 14082 6690
rect 14082 6638 14084 6690
rect 14028 6636 14084 6638
rect 13692 6524 13748 6580
rect 13692 5740 13748 5796
rect 13804 5628 13860 5684
rect 13692 5234 13748 5236
rect 13692 5182 13694 5234
rect 13694 5182 13746 5234
rect 13746 5182 13748 5234
rect 13692 5180 13748 5182
rect 12572 4898 12628 4900
rect 12572 4846 12574 4898
rect 12574 4846 12626 4898
rect 12626 4846 12628 4898
rect 12572 4844 12628 4846
rect 13356 4732 13412 4788
rect 12684 4620 12740 4676
rect 12236 4284 12292 4340
rect 12908 4338 12964 4340
rect 12908 4286 12910 4338
rect 12910 4286 12962 4338
rect 12962 4286 12964 4338
rect 12908 4284 12964 4286
rect 13356 3836 13412 3892
rect 13580 5068 13636 5124
rect 13692 4562 13748 4564
rect 13692 4510 13694 4562
rect 13694 4510 13746 4562
rect 13746 4510 13748 4562
rect 13692 4508 13748 4510
rect 13916 5516 13972 5572
rect 14476 5740 14532 5796
rect 14252 5292 14308 5348
rect 14476 5180 14532 5236
rect 14140 4898 14196 4900
rect 14140 4846 14142 4898
rect 14142 4846 14194 4898
rect 14194 4846 14196 4898
rect 14140 4844 14196 4846
rect 15036 7420 15092 7476
rect 15148 6860 15204 6916
rect 15036 5964 15092 6020
rect 14924 5180 14980 5236
rect 13916 4732 13972 4788
rect 14140 4396 14196 4452
rect 14812 4338 14868 4340
rect 14812 4286 14814 4338
rect 14814 4286 14866 4338
rect 14866 4286 14868 4338
rect 14812 4284 14868 4286
rect 14700 4060 14756 4116
rect 14140 3666 14196 3668
rect 14140 3614 14142 3666
rect 14142 3614 14194 3666
rect 14194 3614 14196 3666
rect 14140 3612 14196 3614
rect 14252 3948 14308 4004
rect 13468 3500 13524 3556
rect 14252 3388 14308 3444
rect 14588 3442 14644 3444
rect 14588 3390 14590 3442
rect 14590 3390 14642 3442
rect 14642 3390 14644 3442
rect 14588 3388 14644 3390
rect 11676 3052 11732 3108
rect 11340 2492 11396 2548
rect 15260 6466 15316 6468
rect 15260 6414 15262 6466
rect 15262 6414 15314 6466
rect 15314 6414 15316 6466
rect 15260 6412 15316 6414
rect 15820 15820 15876 15876
rect 15820 15148 15876 15204
rect 16268 21308 16324 21364
rect 16044 18450 16100 18452
rect 16044 18398 16046 18450
rect 16046 18398 16098 18450
rect 16098 18398 16100 18450
rect 16044 18396 16100 18398
rect 16156 19964 16212 20020
rect 16156 19068 16212 19124
rect 16156 18508 16212 18564
rect 16492 20188 16548 20244
rect 16604 20018 16660 20020
rect 16604 19966 16606 20018
rect 16606 19966 16658 20018
rect 16658 19966 16660 20018
rect 16604 19964 16660 19966
rect 16380 18508 16436 18564
rect 15932 14530 15988 14532
rect 15932 14478 15934 14530
rect 15934 14478 15986 14530
rect 15986 14478 15988 14530
rect 15932 14476 15988 14478
rect 16268 17442 16324 17444
rect 16268 17390 16270 17442
rect 16270 17390 16322 17442
rect 16322 17390 16324 17442
rect 16268 17388 16324 17390
rect 16156 16604 16212 16660
rect 16156 15820 16212 15876
rect 16268 15708 16324 15764
rect 16268 15426 16324 15428
rect 16268 15374 16270 15426
rect 16270 15374 16322 15426
rect 16322 15374 16324 15426
rect 16268 15372 16324 15374
rect 16492 17164 16548 17220
rect 17276 22316 17332 22372
rect 17500 21868 17556 21924
rect 17388 21196 17444 21252
rect 17164 20690 17220 20692
rect 17164 20638 17166 20690
rect 17166 20638 17218 20690
rect 17218 20638 17220 20690
rect 17164 20636 17220 20638
rect 16828 20130 16884 20132
rect 16828 20078 16830 20130
rect 16830 20078 16882 20130
rect 16882 20078 16884 20130
rect 16828 20076 16884 20078
rect 16940 20018 16996 20020
rect 16940 19966 16942 20018
rect 16942 19966 16994 20018
rect 16994 19966 16996 20018
rect 16940 19964 16996 19966
rect 18284 24892 18340 24948
rect 18732 24892 18788 24948
rect 18284 24162 18340 24164
rect 18284 24110 18286 24162
rect 18286 24110 18338 24162
rect 18338 24110 18340 24162
rect 18284 24108 18340 24110
rect 18620 23938 18676 23940
rect 18620 23886 18622 23938
rect 18622 23886 18674 23938
rect 18674 23886 18676 23938
rect 18620 23884 18676 23886
rect 18620 23548 18676 23604
rect 18284 22258 18340 22260
rect 18284 22206 18286 22258
rect 18286 22206 18338 22258
rect 18338 22206 18340 22258
rect 18284 22204 18340 22206
rect 18060 21644 18116 21700
rect 17948 21586 18004 21588
rect 17948 21534 17950 21586
rect 17950 21534 18002 21586
rect 18002 21534 18004 21586
rect 17948 21532 18004 21534
rect 17388 20300 17444 20356
rect 17836 20524 17892 20580
rect 17724 20018 17780 20020
rect 17724 19966 17726 20018
rect 17726 19966 17778 20018
rect 17778 19966 17780 20018
rect 17724 19964 17780 19966
rect 17500 18732 17556 18788
rect 16940 18620 16996 18676
rect 16716 16156 16772 16212
rect 16828 17948 16884 18004
rect 16716 15484 16772 15540
rect 16604 15314 16660 15316
rect 16604 15262 16606 15314
rect 16606 15262 16658 15314
rect 16658 15262 16660 15314
rect 16604 15260 16660 15262
rect 16492 15036 16548 15092
rect 16044 13916 16100 13972
rect 16268 12908 16324 12964
rect 16268 12290 16324 12292
rect 16268 12238 16270 12290
rect 16270 12238 16322 12290
rect 16322 12238 16324 12290
rect 16268 12236 16324 12238
rect 15820 10444 15876 10500
rect 16268 10108 16324 10164
rect 16156 10050 16212 10052
rect 16156 9998 16158 10050
rect 16158 9998 16210 10050
rect 16210 9998 16212 10050
rect 16156 9996 16212 9998
rect 16044 9548 16100 9604
rect 16156 9436 16212 9492
rect 15932 9042 15988 9044
rect 15932 8990 15934 9042
rect 15934 8990 15986 9042
rect 15986 8990 15988 9042
rect 15932 8988 15988 8990
rect 16156 8988 16212 9044
rect 15484 7420 15540 7476
rect 15708 7586 15764 7588
rect 15708 7534 15710 7586
rect 15710 7534 15762 7586
rect 15762 7534 15764 7586
rect 15708 7532 15764 7534
rect 16044 7868 16100 7924
rect 16044 7196 16100 7252
rect 15372 6188 15428 6244
rect 15148 5516 15204 5572
rect 15148 5234 15204 5236
rect 15148 5182 15150 5234
rect 15150 5182 15202 5234
rect 15202 5182 15204 5234
rect 15148 5180 15204 5182
rect 15260 4396 15316 4452
rect 16492 9212 16548 9268
rect 16492 8876 16548 8932
rect 16380 8316 16436 8372
rect 16492 8258 16548 8260
rect 16492 8206 16494 8258
rect 16494 8206 16546 8258
rect 16546 8206 16548 8258
rect 16492 8204 16548 8206
rect 16380 7420 16436 7476
rect 16492 7084 16548 7140
rect 16828 13746 16884 13748
rect 16828 13694 16830 13746
rect 16830 13694 16882 13746
rect 16882 13694 16884 13746
rect 16828 13692 16884 13694
rect 16940 12962 16996 12964
rect 16940 12910 16942 12962
rect 16942 12910 16994 12962
rect 16994 12910 16996 12962
rect 16940 12908 16996 12910
rect 16828 11788 16884 11844
rect 16716 11676 16772 11732
rect 16940 11452 16996 11508
rect 16828 10444 16884 10500
rect 16716 8818 16772 8820
rect 16716 8766 16718 8818
rect 16718 8766 16770 8818
rect 16770 8766 16772 8818
rect 16716 8764 16772 8766
rect 16828 8092 16884 8148
rect 16940 7644 16996 7700
rect 16268 6524 16324 6580
rect 16828 7308 16884 7364
rect 15596 5964 15652 6020
rect 15596 4620 15652 4676
rect 15820 5740 15876 5796
rect 15484 4172 15540 4228
rect 14924 2716 14980 2772
rect 15148 3612 15204 3668
rect 15596 3554 15652 3556
rect 15596 3502 15598 3554
rect 15598 3502 15650 3554
rect 15650 3502 15652 3554
rect 15596 3500 15652 3502
rect 15820 3164 15876 3220
rect 15932 6412 15988 6468
rect 16604 6690 16660 6692
rect 16604 6638 16606 6690
rect 16606 6638 16658 6690
rect 16658 6638 16660 6690
rect 16604 6636 16660 6638
rect 16380 6412 16436 6468
rect 16156 6188 16212 6244
rect 16044 6130 16100 6132
rect 16044 6078 16046 6130
rect 16046 6078 16098 6130
rect 16098 6078 16100 6130
rect 16044 6076 16100 6078
rect 16380 5964 16436 6020
rect 16828 5964 16884 6020
rect 17388 16940 17444 16996
rect 17164 14700 17220 14756
rect 17276 16268 17332 16324
rect 17388 16156 17444 16212
rect 17276 15260 17332 15316
rect 17164 14028 17220 14084
rect 17388 14924 17444 14980
rect 17612 17612 17668 17668
rect 18172 18844 18228 18900
rect 17948 18562 18004 18564
rect 17948 18510 17950 18562
rect 17950 18510 18002 18562
rect 18002 18510 18004 18562
rect 17948 18508 18004 18510
rect 17836 18284 17892 18340
rect 18508 21644 18564 21700
rect 18620 21308 18676 21364
rect 18732 20972 18788 21028
rect 18620 20578 18676 20580
rect 18620 20526 18622 20578
rect 18622 20526 18674 20578
rect 18674 20526 18676 20578
rect 18620 20524 18676 20526
rect 18508 20412 18564 20468
rect 18396 20300 18452 20356
rect 18396 20130 18452 20132
rect 18396 20078 18398 20130
rect 18398 20078 18450 20130
rect 18450 20078 18452 20130
rect 18396 20076 18452 20078
rect 17948 17612 18004 17668
rect 17724 17052 17780 17108
rect 17836 17276 17892 17332
rect 17948 15820 18004 15876
rect 18844 19404 18900 19460
rect 18732 18732 18788 18788
rect 18620 17666 18676 17668
rect 18620 17614 18622 17666
rect 18622 17614 18674 17666
rect 18674 17614 18676 17666
rect 18620 17612 18676 17614
rect 18844 17612 18900 17668
rect 18844 17164 18900 17220
rect 21084 27244 21140 27300
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 25564 19684 25620
rect 19180 24780 19236 24836
rect 20300 25618 20356 25620
rect 20300 25566 20302 25618
rect 20302 25566 20354 25618
rect 20354 25566 20356 25618
rect 20300 25564 20356 25566
rect 20636 25900 20692 25956
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20188 25116 20244 25172
rect 20044 25060 20100 25062
rect 20860 24946 20916 24948
rect 20860 24894 20862 24946
rect 20862 24894 20914 24946
rect 20914 24894 20916 24946
rect 20860 24892 20916 24894
rect 20972 24780 21028 24836
rect 19068 24610 19124 24612
rect 19068 24558 19070 24610
rect 19070 24558 19122 24610
rect 19122 24558 19124 24610
rect 19068 24556 19124 24558
rect 19292 23996 19348 24052
rect 20412 24610 20468 24612
rect 20412 24558 20414 24610
rect 20414 24558 20466 24610
rect 20466 24558 20468 24610
rect 20412 24556 20468 24558
rect 19852 23884 19908 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19068 22316 19124 22372
rect 19292 22204 19348 22260
rect 19404 21644 19460 21700
rect 19180 20524 19236 20580
rect 19180 20188 19236 20244
rect 19068 19628 19124 19684
rect 18956 17276 19012 17332
rect 18284 16828 18340 16884
rect 18172 16156 18228 16212
rect 18284 15820 18340 15876
rect 18508 15596 18564 15652
rect 19068 19404 19124 19460
rect 19292 17948 19348 18004
rect 19180 16604 19236 16660
rect 20300 23154 20356 23156
rect 20300 23102 20302 23154
rect 20302 23102 20354 23154
rect 20354 23102 20356 23154
rect 20300 23100 20356 23102
rect 20972 23660 21028 23716
rect 20076 22652 20132 22708
rect 20524 22316 20580 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 21308 19684 21364
rect 19740 20690 19796 20692
rect 19740 20638 19742 20690
rect 19742 20638 19794 20690
rect 19794 20638 19796 20690
rect 19740 20636 19796 20638
rect 19628 20412 19684 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 19180 20132 19236
rect 19740 19068 19796 19124
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20860 22316 20916 22372
rect 20748 21698 20804 21700
rect 20748 21646 20750 21698
rect 20750 21646 20802 21698
rect 20802 21646 20804 21698
rect 20748 21644 20804 21646
rect 20524 20748 20580 20804
rect 20412 19068 20468 19124
rect 20748 19964 20804 20020
rect 20636 19852 20692 19908
rect 20412 18396 20468 18452
rect 20188 17948 20244 18004
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19852 17052 19908 17108
rect 20076 16322 20132 16324
rect 20076 16270 20078 16322
rect 20078 16270 20130 16322
rect 20130 16270 20132 16322
rect 20076 16268 20132 16270
rect 18844 15932 18900 15988
rect 18732 15090 18788 15092
rect 18732 15038 18734 15090
rect 18734 15038 18786 15090
rect 18786 15038 18788 15090
rect 18732 15036 18788 15038
rect 18396 14700 18452 14756
rect 18172 14588 18228 14644
rect 18396 13916 18452 13972
rect 18732 14700 18788 14756
rect 17612 12348 17668 12404
rect 18060 13746 18116 13748
rect 18060 13694 18062 13746
rect 18062 13694 18114 13746
rect 18114 13694 18116 13746
rect 18060 13692 18116 13694
rect 18172 13580 18228 13636
rect 17836 11676 17892 11732
rect 17612 10892 17668 10948
rect 17724 10834 17780 10836
rect 17724 10782 17726 10834
rect 17726 10782 17778 10834
rect 17778 10782 17780 10834
rect 17724 10780 17780 10782
rect 17388 9826 17444 9828
rect 17388 9774 17390 9826
rect 17390 9774 17442 9826
rect 17442 9774 17444 9826
rect 17388 9772 17444 9774
rect 17164 9436 17220 9492
rect 17164 9100 17220 9156
rect 17500 8316 17556 8372
rect 17276 7756 17332 7812
rect 18060 11170 18116 11172
rect 18060 11118 18062 11170
rect 18062 11118 18114 11170
rect 18114 11118 18116 11170
rect 18060 11116 18116 11118
rect 19964 16098 20020 16100
rect 19964 16046 19966 16098
rect 19966 16046 20018 16098
rect 20018 16046 20020 16098
rect 19964 16044 20020 16046
rect 19628 15820 19684 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18956 15372 19012 15428
rect 18732 13356 18788 13412
rect 18284 12348 18340 12404
rect 18620 11228 18676 11284
rect 18620 10892 18676 10948
rect 17948 10610 18004 10612
rect 17948 10558 17950 10610
rect 17950 10558 18002 10610
rect 18002 10558 18004 10610
rect 17948 10556 18004 10558
rect 18060 10498 18116 10500
rect 18060 10446 18062 10498
rect 18062 10446 18114 10498
rect 18114 10446 18116 10498
rect 18060 10444 18116 10446
rect 17836 9154 17892 9156
rect 17836 9102 17838 9154
rect 17838 9102 17890 9154
rect 17890 9102 17892 9154
rect 17836 9100 17892 9102
rect 18172 9714 18228 9716
rect 18172 9662 18174 9714
rect 18174 9662 18226 9714
rect 18226 9662 18228 9714
rect 18172 9660 18228 9662
rect 18060 8818 18116 8820
rect 18060 8766 18062 8818
rect 18062 8766 18114 8818
rect 18114 8766 18116 8818
rect 18060 8764 18116 8766
rect 18172 8652 18228 8708
rect 16492 5292 16548 5348
rect 16716 5234 16772 5236
rect 16716 5182 16718 5234
rect 16718 5182 16770 5234
rect 16770 5182 16772 5234
rect 16716 5180 16772 5182
rect 16044 4562 16100 4564
rect 16044 4510 16046 4562
rect 16046 4510 16098 4562
rect 16098 4510 16100 4562
rect 16044 4508 16100 4510
rect 16940 5346 16996 5348
rect 16940 5294 16942 5346
rect 16942 5294 16994 5346
rect 16994 5294 16996 5346
rect 16940 5292 16996 5294
rect 16604 4508 16660 4564
rect 16268 4338 16324 4340
rect 16268 4286 16270 4338
rect 16270 4286 16322 4338
rect 16322 4286 16324 4338
rect 16268 4284 16324 4286
rect 16492 3836 16548 3892
rect 16044 3666 16100 3668
rect 16044 3614 16046 3666
rect 16046 3614 16098 3666
rect 16098 3614 16100 3666
rect 16044 3612 16100 3614
rect 17276 5964 17332 6020
rect 17052 3724 17108 3780
rect 17164 4284 17220 4340
rect 17500 6860 17556 6916
rect 17500 5852 17556 5908
rect 17836 7980 17892 8036
rect 17948 8204 18004 8260
rect 18620 10220 18676 10276
rect 18396 9436 18452 9492
rect 18620 9660 18676 9716
rect 18508 8204 18564 8260
rect 19404 15036 19460 15092
rect 19292 14588 19348 14644
rect 19068 12684 19124 12740
rect 19068 12460 19124 12516
rect 19180 12124 19236 12180
rect 18956 11676 19012 11732
rect 19068 11506 19124 11508
rect 19068 11454 19070 11506
rect 19070 11454 19122 11506
rect 19122 11454 19124 11506
rect 19068 11452 19124 11454
rect 18844 11340 18900 11396
rect 19964 15314 20020 15316
rect 19964 15262 19966 15314
rect 19966 15262 20018 15314
rect 20018 15262 20020 15314
rect 19964 15260 20020 15262
rect 19852 15036 19908 15092
rect 20524 18284 20580 18340
rect 20748 19010 20804 19012
rect 20748 18958 20750 19010
rect 20750 18958 20802 19010
rect 20802 18958 20804 19010
rect 20748 18956 20804 18958
rect 20748 18450 20804 18452
rect 20748 18398 20750 18450
rect 20750 18398 20802 18450
rect 20802 18398 20804 18450
rect 20748 18396 20804 18398
rect 20636 17836 20692 17892
rect 20300 17276 20356 17332
rect 20300 16882 20356 16884
rect 20300 16830 20302 16882
rect 20302 16830 20354 16882
rect 20354 16830 20356 16882
rect 20300 16828 20356 16830
rect 20748 17164 20804 17220
rect 20524 16380 20580 16436
rect 21644 26572 21700 26628
rect 21196 26402 21252 26404
rect 21196 26350 21198 26402
rect 21198 26350 21250 26402
rect 21250 26350 21252 26402
rect 21196 26348 21252 26350
rect 22764 27074 22820 27076
rect 22764 27022 22766 27074
rect 22766 27022 22818 27074
rect 22818 27022 22820 27074
rect 22764 27020 22820 27022
rect 22876 26850 22932 26852
rect 22876 26798 22878 26850
rect 22878 26798 22930 26850
rect 22930 26798 22932 26850
rect 22876 26796 22932 26798
rect 24220 27746 24276 27748
rect 24220 27694 24222 27746
rect 24222 27694 24274 27746
rect 24274 27694 24276 27746
rect 24220 27692 24276 27694
rect 25228 27692 25284 27748
rect 29596 31612 29652 31668
rect 26684 29986 26740 29988
rect 26684 29934 26686 29986
rect 26686 29934 26738 29986
rect 26738 29934 26740 29986
rect 26684 29932 26740 29934
rect 27916 29314 27972 29316
rect 27916 29262 27918 29314
rect 27918 29262 27970 29314
rect 27970 29262 27972 29314
rect 27916 29260 27972 29262
rect 28364 29260 28420 29316
rect 28588 29650 28644 29652
rect 28588 29598 28590 29650
rect 28590 29598 28642 29650
rect 28642 29598 28644 29650
rect 28588 29596 28644 29598
rect 26572 28588 26628 28644
rect 27916 28588 27972 28644
rect 27692 28530 27748 28532
rect 27692 28478 27694 28530
rect 27694 28478 27746 28530
rect 27746 28478 27748 28530
rect 27692 28476 27748 28478
rect 26124 28364 26180 28420
rect 26012 28082 26068 28084
rect 26012 28030 26014 28082
rect 26014 28030 26066 28082
rect 26066 28030 26068 28082
rect 26012 28028 26068 28030
rect 26684 28028 26740 28084
rect 21756 26236 21812 26292
rect 22092 26012 22148 26068
rect 21420 25900 21476 25956
rect 22540 25730 22596 25732
rect 22540 25678 22542 25730
rect 22542 25678 22594 25730
rect 22594 25678 22596 25730
rect 22540 25676 22596 25678
rect 23436 26572 23492 26628
rect 23548 26796 23604 26852
rect 22876 26124 22932 26180
rect 22988 25788 23044 25844
rect 22764 25564 22820 25620
rect 23436 26012 23492 26068
rect 23100 25618 23156 25620
rect 23100 25566 23102 25618
rect 23102 25566 23154 25618
rect 23154 25566 23156 25618
rect 23100 25564 23156 25566
rect 23324 25004 23380 25060
rect 22876 24444 22932 24500
rect 24332 26796 24388 26852
rect 24220 26290 24276 26292
rect 24220 26238 24222 26290
rect 24222 26238 24274 26290
rect 24274 26238 24276 26290
rect 24220 26236 24276 26238
rect 24780 26572 24836 26628
rect 23996 26178 24052 26180
rect 23996 26126 23998 26178
rect 23998 26126 24050 26178
rect 24050 26126 24052 26178
rect 23996 26124 24052 26126
rect 23772 25788 23828 25844
rect 23884 25676 23940 25732
rect 24668 25618 24724 25620
rect 24668 25566 24670 25618
rect 24670 25566 24722 25618
rect 24722 25566 24724 25618
rect 24668 25564 24724 25566
rect 25900 26124 25956 26180
rect 27132 28028 27188 28084
rect 29148 28642 29204 28644
rect 29148 28590 29150 28642
rect 29150 28590 29202 28642
rect 29202 28590 29204 28642
rect 29148 28588 29204 28590
rect 28140 28476 28196 28532
rect 30156 30940 30212 30996
rect 29372 28476 29428 28532
rect 29484 28588 29540 28644
rect 32396 35026 32452 35028
rect 32396 34974 32398 35026
rect 32398 34974 32450 35026
rect 32450 34974 32452 35026
rect 32396 34972 32452 34974
rect 34300 38108 34356 38164
rect 34524 38050 34580 38052
rect 34524 37998 34526 38050
rect 34526 37998 34578 38050
rect 34578 37998 34580 38050
rect 34524 37996 34580 37998
rect 34636 37938 34692 37940
rect 34636 37886 34638 37938
rect 34638 37886 34690 37938
rect 34690 37886 34692 37938
rect 34636 37884 34692 37886
rect 34300 37548 34356 37604
rect 34188 37100 34244 37156
rect 34412 37266 34468 37268
rect 34412 37214 34414 37266
rect 34414 37214 34466 37266
rect 34466 37214 34468 37266
rect 34412 37212 34468 37214
rect 34748 37154 34804 37156
rect 34748 37102 34750 37154
rect 34750 37102 34802 37154
rect 34802 37102 34804 37154
rect 34748 37100 34804 37102
rect 36876 39788 36932 39844
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 38050 35140 38052
rect 35084 37998 35086 38050
rect 35086 37998 35138 38050
rect 35138 37998 35140 38050
rect 35084 37996 35140 37998
rect 35196 37266 35252 37268
rect 35196 37214 35198 37266
rect 35198 37214 35250 37266
rect 35250 37214 35252 37266
rect 35196 37212 35252 37214
rect 35644 37772 35700 37828
rect 35420 37100 35476 37156
rect 35756 37100 35812 37156
rect 34972 37042 35028 37044
rect 34972 36990 34974 37042
rect 34974 36990 35026 37042
rect 35026 36990 35028 37042
rect 34972 36988 35028 36990
rect 34636 36428 34692 36484
rect 34188 35980 34244 36036
rect 34524 35868 34580 35924
rect 34636 35420 34692 35476
rect 32508 34802 32564 34804
rect 32508 34750 32510 34802
rect 32510 34750 32562 34802
rect 32562 34750 32564 34802
rect 32508 34748 32564 34750
rect 34636 34636 34692 34692
rect 33404 34354 33460 34356
rect 33404 34302 33406 34354
rect 33406 34302 33458 34354
rect 33458 34302 33460 34354
rect 33404 34300 33460 34302
rect 33852 34354 33908 34356
rect 33852 34302 33854 34354
rect 33854 34302 33906 34354
rect 33906 34302 33908 34354
rect 33852 34300 33908 34302
rect 32172 34130 32228 34132
rect 32172 34078 32174 34130
rect 32174 34078 32226 34130
rect 32226 34078 32228 34130
rect 32172 34076 32228 34078
rect 32172 33346 32228 33348
rect 32172 33294 32174 33346
rect 32174 33294 32226 33346
rect 32226 33294 32228 33346
rect 32172 33292 32228 33294
rect 34412 34130 34468 34132
rect 34412 34078 34414 34130
rect 34414 34078 34466 34130
rect 34466 34078 34468 34130
rect 34412 34076 34468 34078
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35644 36482 35700 36484
rect 35644 36430 35646 36482
rect 35646 36430 35698 36482
rect 35698 36430 35700 36482
rect 35644 36428 35700 36430
rect 35532 36316 35588 36372
rect 34860 35922 34916 35924
rect 34860 35870 34862 35922
rect 34862 35870 34914 35922
rect 34914 35870 34916 35922
rect 34860 35868 34916 35870
rect 35644 35922 35700 35924
rect 35644 35870 35646 35922
rect 35646 35870 35698 35922
rect 35698 35870 35700 35922
rect 35644 35868 35700 35870
rect 34972 35756 35028 35812
rect 36204 35868 36260 35924
rect 36428 35756 36484 35812
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34972 35084 35028 35140
rect 34860 34690 34916 34692
rect 34860 34638 34862 34690
rect 34862 34638 34914 34690
rect 34914 34638 34916 34690
rect 34860 34636 34916 34638
rect 35084 34914 35140 34916
rect 35084 34862 35086 34914
rect 35086 34862 35138 34914
rect 35138 34862 35140 34914
rect 35084 34860 35140 34862
rect 37324 42924 37380 42980
rect 37548 43372 37604 43428
rect 38556 48354 38612 48356
rect 38556 48302 38558 48354
rect 38558 48302 38610 48354
rect 38610 48302 38612 48354
rect 38556 48300 38612 48302
rect 38332 48242 38388 48244
rect 38332 48190 38334 48242
rect 38334 48190 38386 48242
rect 38386 48190 38388 48242
rect 38332 48188 38388 48190
rect 38108 47346 38164 47348
rect 38108 47294 38110 47346
rect 38110 47294 38162 47346
rect 38162 47294 38164 47346
rect 38108 47292 38164 47294
rect 39116 48242 39172 48244
rect 39116 48190 39118 48242
rect 39118 48190 39170 48242
rect 39170 48190 39172 48242
rect 39116 48188 39172 48190
rect 39900 50482 39956 50484
rect 39900 50430 39902 50482
rect 39902 50430 39954 50482
rect 39954 50430 39956 50482
rect 39900 50428 39956 50430
rect 39564 49138 39620 49140
rect 39564 49086 39566 49138
rect 39566 49086 39618 49138
rect 39618 49086 39620 49138
rect 39564 49084 39620 49086
rect 39452 49026 39508 49028
rect 39452 48974 39454 49026
rect 39454 48974 39506 49026
rect 39506 48974 39508 49026
rect 39452 48972 39508 48974
rect 39452 48242 39508 48244
rect 39452 48190 39454 48242
rect 39454 48190 39506 48242
rect 39506 48190 39508 48242
rect 39452 48188 39508 48190
rect 40908 51154 40964 51156
rect 40908 51102 40910 51154
rect 40910 51102 40962 51154
rect 40962 51102 40964 51154
rect 40908 51100 40964 51102
rect 41132 51324 41188 51380
rect 42252 52162 42308 52164
rect 42252 52110 42254 52162
rect 42254 52110 42306 52162
rect 42306 52110 42308 52162
rect 42252 52108 42308 52110
rect 42028 51436 42084 51492
rect 42140 51660 42196 51716
rect 39788 48300 39844 48356
rect 40236 48524 40292 48580
rect 40012 48188 40068 48244
rect 40236 48076 40292 48132
rect 39340 47180 39396 47236
rect 39116 47068 39172 47124
rect 40124 47964 40180 48020
rect 41020 48130 41076 48132
rect 41020 48078 41022 48130
rect 41022 48078 41074 48130
rect 41074 48078 41076 48130
rect 41020 48076 41076 48078
rect 40236 47516 40292 47572
rect 39900 46844 39956 46900
rect 40012 47068 40068 47124
rect 37996 45218 38052 45220
rect 37996 45166 37998 45218
rect 37998 45166 38050 45218
rect 38050 45166 38052 45218
rect 37996 45164 38052 45166
rect 37884 45106 37940 45108
rect 37884 45054 37886 45106
rect 37886 45054 37938 45106
rect 37938 45054 37940 45106
rect 37884 45052 37940 45054
rect 38780 44716 38836 44772
rect 39452 45778 39508 45780
rect 39452 45726 39454 45778
rect 39454 45726 39506 45778
rect 39506 45726 39508 45778
rect 39452 45724 39508 45726
rect 41020 46898 41076 46900
rect 41020 46846 41022 46898
rect 41022 46846 41074 46898
rect 41074 46846 41076 46898
rect 41020 46844 41076 46846
rect 39452 45106 39508 45108
rect 39452 45054 39454 45106
rect 39454 45054 39506 45106
rect 39506 45054 39508 45106
rect 39452 45052 39508 45054
rect 39116 44828 39172 44884
rect 38668 44380 38724 44436
rect 39788 44940 39844 44996
rect 39676 44434 39732 44436
rect 39676 44382 39678 44434
rect 39678 44382 39730 44434
rect 39730 44382 39732 44434
rect 39676 44380 39732 44382
rect 38332 43820 38388 43876
rect 38108 43538 38164 43540
rect 38108 43486 38110 43538
rect 38110 43486 38162 43538
rect 38162 43486 38164 43538
rect 38108 43484 38164 43486
rect 37884 43426 37940 43428
rect 37884 43374 37886 43426
rect 37886 43374 37938 43426
rect 37938 43374 37940 43426
rect 37884 43372 37940 43374
rect 37884 42924 37940 42980
rect 37212 39452 37268 39508
rect 37436 39506 37492 39508
rect 37436 39454 37438 39506
rect 37438 39454 37490 39506
rect 37490 39454 37492 39506
rect 37436 39452 37492 39454
rect 38780 44268 38836 44324
rect 39228 44210 39284 44212
rect 39228 44158 39230 44210
rect 39230 44158 39282 44210
rect 39282 44158 39284 44210
rect 39228 44156 39284 44158
rect 44828 55186 44884 55188
rect 44828 55134 44830 55186
rect 44830 55134 44882 55186
rect 44882 55134 44884 55186
rect 44828 55132 44884 55134
rect 44940 55074 44996 55076
rect 44940 55022 44942 55074
rect 44942 55022 44994 55074
rect 44994 55022 44996 55074
rect 44940 55020 44996 55022
rect 45164 55074 45220 55076
rect 45164 55022 45166 55074
rect 45166 55022 45218 55074
rect 45218 55022 45220 55074
rect 45164 55020 45220 55022
rect 45500 55186 45556 55188
rect 45500 55134 45502 55186
rect 45502 55134 45554 55186
rect 45554 55134 45556 55186
rect 45500 55132 45556 55134
rect 45724 55186 45780 55188
rect 45724 55134 45726 55186
rect 45726 55134 45778 55186
rect 45778 55134 45780 55186
rect 45724 55132 45780 55134
rect 43484 54514 43540 54516
rect 43484 54462 43486 54514
rect 43486 54462 43538 54514
rect 43538 54462 43540 54514
rect 43484 54460 43540 54462
rect 43596 53788 43652 53844
rect 44380 54514 44436 54516
rect 44380 54462 44382 54514
rect 44382 54462 44434 54514
rect 44434 54462 44436 54514
rect 44380 54460 44436 54462
rect 43820 53788 43876 53844
rect 43932 53618 43988 53620
rect 43932 53566 43934 53618
rect 43934 53566 43986 53618
rect 43986 53566 43988 53618
rect 43932 53564 43988 53566
rect 46844 54626 46900 54628
rect 46844 54574 46846 54626
rect 46846 54574 46898 54626
rect 46898 54574 46900 54626
rect 46844 54572 46900 54574
rect 46172 53954 46228 53956
rect 46172 53902 46174 53954
rect 46174 53902 46226 53954
rect 46226 53902 46228 53954
rect 46172 53900 46228 53902
rect 44828 53564 44884 53620
rect 47068 55186 47124 55188
rect 47068 55134 47070 55186
rect 47070 55134 47122 55186
rect 47122 55134 47124 55186
rect 47068 55132 47124 55134
rect 46956 54124 47012 54180
rect 47628 54572 47684 54628
rect 47516 54124 47572 54180
rect 42588 52108 42644 52164
rect 43148 51660 43204 51716
rect 42476 50594 42532 50596
rect 42476 50542 42478 50594
rect 42478 50542 42530 50594
rect 42530 50542 42532 50594
rect 42476 50540 42532 50542
rect 43484 50540 43540 50596
rect 43932 52108 43988 52164
rect 44940 52108 44996 52164
rect 44044 51266 44100 51268
rect 44044 51214 44046 51266
rect 44046 51214 44098 51266
rect 44098 51214 44100 51266
rect 44044 51212 44100 51214
rect 44268 50876 44324 50932
rect 44156 50482 44212 50484
rect 44156 50430 44158 50482
rect 44158 50430 44210 50482
rect 44210 50430 44212 50482
rect 44156 50428 44212 50430
rect 43036 49922 43092 49924
rect 43036 49870 43038 49922
rect 43038 49870 43090 49922
rect 43090 49870 43092 49922
rect 43036 49868 43092 49870
rect 43372 49810 43428 49812
rect 43372 49758 43374 49810
rect 43374 49758 43426 49810
rect 43426 49758 43428 49810
rect 43372 49756 43428 49758
rect 42252 49026 42308 49028
rect 42252 48974 42254 49026
rect 42254 48974 42306 49026
rect 42306 48974 42308 49026
rect 42252 48972 42308 48974
rect 42812 49026 42868 49028
rect 42812 48974 42814 49026
rect 42814 48974 42866 49026
rect 42866 48974 42868 49026
rect 42812 48972 42868 48974
rect 43260 49026 43316 49028
rect 43260 48974 43262 49026
rect 43262 48974 43314 49026
rect 43314 48974 43316 49026
rect 43260 48972 43316 48974
rect 42924 48914 42980 48916
rect 42924 48862 42926 48914
rect 42926 48862 42978 48914
rect 42978 48862 42980 48914
rect 42924 48860 42980 48862
rect 43036 48748 43092 48804
rect 42140 48354 42196 48356
rect 42140 48302 42142 48354
rect 42142 48302 42194 48354
rect 42194 48302 42196 48354
rect 42140 48300 42196 48302
rect 42476 48354 42532 48356
rect 42476 48302 42478 48354
rect 42478 48302 42530 48354
rect 42530 48302 42532 48354
rect 42476 48300 42532 48302
rect 42028 46786 42084 46788
rect 42028 46734 42030 46786
rect 42030 46734 42082 46786
rect 42082 46734 42084 46786
rect 42028 46732 42084 46734
rect 41244 45276 41300 45332
rect 40460 44380 40516 44436
rect 40908 45164 40964 45220
rect 40124 44156 40180 44212
rect 38668 42924 38724 42980
rect 38556 42754 38612 42756
rect 38556 42702 38558 42754
rect 38558 42702 38610 42754
rect 38610 42702 38612 42754
rect 38556 42700 38612 42702
rect 38668 42194 38724 42196
rect 38668 42142 38670 42194
rect 38670 42142 38722 42194
rect 38722 42142 38724 42194
rect 38668 42140 38724 42142
rect 39228 43260 39284 43316
rect 39004 42754 39060 42756
rect 39004 42702 39006 42754
rect 39006 42702 39058 42754
rect 39058 42702 39060 42754
rect 39004 42700 39060 42702
rect 39900 42754 39956 42756
rect 39900 42702 39902 42754
rect 39902 42702 39954 42754
rect 39954 42702 39956 42754
rect 39900 42700 39956 42702
rect 38444 39788 38500 39844
rect 37996 38556 38052 38612
rect 36988 37548 37044 37604
rect 37212 37826 37268 37828
rect 37212 37774 37214 37826
rect 37214 37774 37266 37826
rect 37266 37774 37268 37826
rect 37212 37772 37268 37774
rect 36876 36876 36932 36932
rect 36876 36428 36932 36484
rect 35980 35084 36036 35140
rect 35868 34914 35924 34916
rect 35868 34862 35870 34914
rect 35870 34862 35922 34914
rect 35922 34862 35924 34914
rect 35868 34860 35924 34862
rect 36988 34076 37044 34132
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 33068 33292 33124 33348
rect 35644 33346 35700 33348
rect 35644 33294 35646 33346
rect 35646 33294 35698 33346
rect 35698 33294 35700 33346
rect 35644 33292 35700 33294
rect 37884 36652 37940 36708
rect 37884 36482 37940 36484
rect 37884 36430 37886 36482
rect 37886 36430 37938 36482
rect 37938 36430 37940 36482
rect 37884 36428 37940 36430
rect 37996 36370 38052 36372
rect 37996 36318 37998 36370
rect 37998 36318 38050 36370
rect 38050 36318 38052 36370
rect 37996 36316 38052 36318
rect 37996 36092 38052 36148
rect 31500 30940 31556 30996
rect 31612 32674 31668 32676
rect 31612 32622 31614 32674
rect 31614 32622 31666 32674
rect 31666 32622 31668 32674
rect 31612 32620 31668 32622
rect 32956 30994 33012 30996
rect 32956 30942 32958 30994
rect 32958 30942 33010 30994
rect 33010 30942 33012 30994
rect 32956 30940 33012 30942
rect 31612 30044 31668 30100
rect 33068 30380 33124 30436
rect 31276 29372 31332 29428
rect 30268 28588 30324 28644
rect 32732 28530 32788 28532
rect 32732 28478 32734 28530
rect 32734 28478 32786 28530
rect 32786 28478 32788 28530
rect 32732 28476 32788 28478
rect 26908 27468 26964 27524
rect 24780 25452 24836 25508
rect 25340 26066 25396 26068
rect 25340 26014 25342 26066
rect 25342 26014 25394 26066
rect 25394 26014 25396 26066
rect 25340 26012 25396 26014
rect 26124 26012 26180 26068
rect 26684 26124 26740 26180
rect 25788 25340 25844 25396
rect 23884 25116 23940 25172
rect 23324 24498 23380 24500
rect 23324 24446 23326 24498
rect 23326 24446 23378 24498
rect 23378 24446 23380 24498
rect 23324 24444 23380 24446
rect 23548 24498 23604 24500
rect 23548 24446 23550 24498
rect 23550 24446 23602 24498
rect 23602 24446 23604 24498
rect 23548 24444 23604 24446
rect 22876 24108 22932 24164
rect 23324 24108 23380 24164
rect 21420 23996 21476 24052
rect 22988 23938 23044 23940
rect 22988 23886 22990 23938
rect 22990 23886 23042 23938
rect 23042 23886 23044 23938
rect 22988 23884 23044 23886
rect 22876 23826 22932 23828
rect 22876 23774 22878 23826
rect 22878 23774 22930 23826
rect 22930 23774 22932 23826
rect 22876 23772 22932 23774
rect 21420 23100 21476 23156
rect 21980 23548 22036 23604
rect 21532 22316 21588 22372
rect 21644 21756 21700 21812
rect 21980 22428 22036 22484
rect 22428 21868 22484 21924
rect 22540 22988 22596 23044
rect 22316 21756 22372 21812
rect 21868 21644 21924 21700
rect 22428 20972 22484 21028
rect 21532 20690 21588 20692
rect 21532 20638 21534 20690
rect 21534 20638 21586 20690
rect 21586 20638 21588 20690
rect 21532 20636 21588 20638
rect 21420 20412 21476 20468
rect 21756 20300 21812 20356
rect 21308 20076 21364 20132
rect 21532 20018 21588 20020
rect 21532 19966 21534 20018
rect 21534 19966 21586 20018
rect 21586 19966 21588 20018
rect 21532 19964 21588 19966
rect 21308 19628 21364 19684
rect 21532 19292 21588 19348
rect 22092 19516 22148 19572
rect 21756 18956 21812 19012
rect 21308 18508 21364 18564
rect 21980 18396 22036 18452
rect 21756 18172 21812 18228
rect 21532 17948 21588 18004
rect 20860 16380 20916 16436
rect 21196 17164 21252 17220
rect 20972 16268 21028 16324
rect 20188 14812 20244 14868
rect 19852 14700 19908 14756
rect 19740 14252 19796 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19292 11452 19348 11508
rect 19404 13580 19460 13636
rect 19068 10892 19124 10948
rect 19180 10668 19236 10724
rect 19292 10556 19348 10612
rect 19068 10220 19124 10276
rect 19068 9100 19124 9156
rect 19852 13804 19908 13860
rect 19852 13020 19908 13076
rect 21308 15874 21364 15876
rect 21308 15822 21310 15874
rect 21310 15822 21362 15874
rect 21362 15822 21364 15874
rect 21308 15820 21364 15822
rect 23100 23714 23156 23716
rect 23100 23662 23102 23714
rect 23102 23662 23154 23714
rect 23154 23662 23156 23714
rect 23100 23660 23156 23662
rect 25004 24668 25060 24724
rect 26012 24722 26068 24724
rect 26012 24670 26014 24722
rect 26014 24670 26066 24722
rect 26066 24670 26068 24722
rect 26012 24668 26068 24670
rect 24556 24444 24612 24500
rect 23772 23826 23828 23828
rect 23772 23774 23774 23826
rect 23774 23774 23826 23826
rect 23826 23774 23828 23826
rect 23772 23772 23828 23774
rect 22764 21756 22820 21812
rect 22988 21810 23044 21812
rect 22988 21758 22990 21810
rect 22990 21758 23042 21810
rect 23042 21758 23044 21810
rect 22988 21756 23044 21758
rect 22652 21196 22708 21252
rect 23100 21196 23156 21252
rect 22876 20972 22932 21028
rect 22316 20412 22372 20468
rect 23324 20412 23380 20468
rect 23212 20188 23268 20244
rect 22428 19292 22484 19348
rect 21868 17388 21924 17444
rect 21420 15314 21476 15316
rect 21420 15262 21422 15314
rect 21422 15262 21474 15314
rect 21474 15262 21476 15314
rect 21420 15260 21476 15262
rect 20188 12684 20244 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19852 12236 19908 12292
rect 20076 11788 20132 11844
rect 19852 11452 19908 11508
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19740 10332 19796 10388
rect 20188 10444 20244 10500
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 8818 19572 8820
rect 19516 8766 19518 8818
rect 19518 8766 19570 8818
rect 19570 8766 19572 8818
rect 19516 8764 19572 8766
rect 18844 8204 18900 8260
rect 17836 7308 17892 7364
rect 18508 7362 18564 7364
rect 18508 7310 18510 7362
rect 18510 7310 18562 7362
rect 18562 7310 18564 7362
rect 18508 7308 18564 7310
rect 18732 7250 18788 7252
rect 18732 7198 18734 7250
rect 18734 7198 18786 7250
rect 18786 7198 18788 7250
rect 18732 7196 18788 7198
rect 18396 6690 18452 6692
rect 18396 6638 18398 6690
rect 18398 6638 18450 6690
rect 18450 6638 18452 6690
rect 18396 6636 18452 6638
rect 18060 6018 18116 6020
rect 18060 5966 18062 6018
rect 18062 5966 18114 6018
rect 18114 5966 18116 6018
rect 18060 5964 18116 5966
rect 18284 6524 18340 6580
rect 17724 4562 17780 4564
rect 17724 4510 17726 4562
rect 17726 4510 17778 4562
rect 17778 4510 17780 4562
rect 17724 4508 17780 4510
rect 17724 3666 17780 3668
rect 17724 3614 17726 3666
rect 17726 3614 17778 3666
rect 17778 3614 17780 3666
rect 17724 3612 17780 3614
rect 17276 3052 17332 3108
rect 15932 2940 15988 2996
rect 15372 2828 15428 2884
rect 15148 2716 15204 2772
rect 17948 5404 18004 5460
rect 18396 5628 18452 5684
rect 18620 5516 18676 5572
rect 18284 5122 18340 5124
rect 18284 5070 18286 5122
rect 18286 5070 18338 5122
rect 18338 5070 18340 5122
rect 18284 5068 18340 5070
rect 18060 4898 18116 4900
rect 18060 4846 18062 4898
rect 18062 4846 18114 4898
rect 18114 4846 18116 4898
rect 18060 4844 18116 4846
rect 18284 4732 18340 4788
rect 17836 3164 17892 3220
rect 17724 2604 17780 2660
rect 18396 3612 18452 3668
rect 18508 4508 18564 4564
rect 20636 12962 20692 12964
rect 20636 12910 20638 12962
rect 20638 12910 20690 12962
rect 20690 12910 20692 12962
rect 20636 12908 20692 12910
rect 20412 11788 20468 11844
rect 20524 12572 20580 12628
rect 20748 12178 20804 12180
rect 20748 12126 20750 12178
rect 20750 12126 20802 12178
rect 20802 12126 20804 12178
rect 20748 12124 20804 12126
rect 21308 14700 21364 14756
rect 21532 14812 21588 14868
rect 21196 13634 21252 13636
rect 21196 13582 21198 13634
rect 21198 13582 21250 13634
rect 21250 13582 21252 13634
rect 21196 13580 21252 13582
rect 21196 13020 21252 13076
rect 20524 10780 20580 10836
rect 20636 11788 20692 11844
rect 20412 10556 20468 10612
rect 20524 9996 20580 10052
rect 21420 12236 21476 12292
rect 20748 10892 20804 10948
rect 20860 9884 20916 9940
rect 20524 8652 20580 8708
rect 20412 8540 20468 8596
rect 19292 8204 19348 8260
rect 20188 8146 20244 8148
rect 20188 8094 20190 8146
rect 20190 8094 20242 8146
rect 20242 8094 20244 8146
rect 20188 8092 20244 8094
rect 19516 7980 19572 8036
rect 19068 7868 19124 7924
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20300 7868 20356 7924
rect 19180 7196 19236 7252
rect 18956 7084 19012 7140
rect 18956 6300 19012 6356
rect 19180 6972 19236 7028
rect 20300 7420 20356 7476
rect 19852 6860 19908 6916
rect 19964 6636 20020 6692
rect 20188 6972 20244 7028
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18844 5628 18900 5684
rect 19180 6018 19236 6020
rect 19180 5966 19182 6018
rect 19182 5966 19234 6018
rect 19234 5966 19236 6018
rect 19180 5964 19236 5966
rect 19068 5740 19124 5796
rect 19068 5516 19124 5572
rect 19404 6130 19460 6132
rect 19404 6078 19406 6130
rect 19406 6078 19458 6130
rect 19458 6078 19460 6130
rect 19404 6076 19460 6078
rect 19292 4844 19348 4900
rect 18956 4226 19012 4228
rect 18956 4174 18958 4226
rect 18958 4174 19010 4226
rect 19010 4174 19012 4226
rect 18956 4172 19012 4174
rect 18956 3666 19012 3668
rect 18956 3614 18958 3666
rect 18958 3614 19010 3666
rect 19010 3614 19012 3666
rect 18956 3612 19012 3614
rect 18060 2492 18116 2548
rect 14924 2156 14980 2212
rect 19292 4338 19348 4340
rect 19292 4286 19294 4338
rect 19294 4286 19346 4338
rect 19346 4286 19348 4338
rect 19292 4284 19348 4286
rect 19180 3948 19236 4004
rect 19628 5292 19684 5348
rect 20524 7586 20580 7588
rect 20524 7534 20526 7586
rect 20526 7534 20578 7586
rect 20578 7534 20580 7586
rect 20524 7532 20580 7534
rect 20636 7420 20692 7476
rect 20412 5516 20468 5572
rect 19516 4732 19572 4788
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19964 4338 20020 4340
rect 19964 4286 19966 4338
rect 19966 4286 20018 4338
rect 20018 4286 20020 4338
rect 19964 4284 20020 4286
rect 20300 3724 20356 3780
rect 19180 3500 19236 3556
rect 19852 3442 19908 3444
rect 19852 3390 19854 3442
rect 19854 3390 19906 3442
rect 19906 3390 19908 3442
rect 19852 3388 19908 3390
rect 20636 5852 20692 5908
rect 21308 10220 21364 10276
rect 21084 9772 21140 9828
rect 21084 8428 21140 8484
rect 21196 9436 21252 9492
rect 21084 8092 21140 8148
rect 21084 7196 21140 7252
rect 21868 12962 21924 12964
rect 21868 12910 21870 12962
rect 21870 12910 21922 12962
rect 21922 12910 21924 12962
rect 21868 12908 21924 12910
rect 22204 16716 22260 16772
rect 22540 18172 22596 18228
rect 22540 17052 22596 17108
rect 22092 15986 22148 15988
rect 22092 15934 22094 15986
rect 22094 15934 22146 15986
rect 22146 15934 22148 15986
rect 22092 15932 22148 15934
rect 22316 15820 22372 15876
rect 22316 15596 22372 15652
rect 22092 12124 22148 12180
rect 21980 11900 22036 11956
rect 21868 11788 21924 11844
rect 21644 11452 21700 11508
rect 22316 12012 22372 12068
rect 21756 9826 21812 9828
rect 21756 9774 21758 9826
rect 21758 9774 21810 9826
rect 21810 9774 21812 9826
rect 21756 9772 21812 9774
rect 21532 8988 21588 9044
rect 21420 8204 21476 8260
rect 21644 8146 21700 8148
rect 21644 8094 21646 8146
rect 21646 8094 21698 8146
rect 21698 8094 21700 8146
rect 21644 8092 21700 8094
rect 20860 5628 20916 5684
rect 21308 6972 21364 7028
rect 20860 4732 20916 4788
rect 20972 4844 21028 4900
rect 21196 6748 21252 6804
rect 21308 6636 21364 6692
rect 21420 6412 21476 6468
rect 21308 5404 21364 5460
rect 21420 6188 21476 6244
rect 21532 5740 21588 5796
rect 21196 5180 21252 5236
rect 21308 5122 21364 5124
rect 21308 5070 21310 5122
rect 21310 5070 21362 5122
rect 21362 5070 21364 5122
rect 21308 5068 21364 5070
rect 20972 3836 21028 3892
rect 21420 4396 21476 4452
rect 21420 3836 21476 3892
rect 21868 8876 21924 8932
rect 22204 10610 22260 10612
rect 22204 10558 22206 10610
rect 22206 10558 22258 10610
rect 22258 10558 22260 10610
rect 22204 10556 22260 10558
rect 22540 16716 22596 16772
rect 22540 15708 22596 15764
rect 22764 19516 22820 19572
rect 22988 17276 23044 17332
rect 22652 16156 22708 16212
rect 22764 16044 22820 16100
rect 22652 15596 22708 15652
rect 22764 15314 22820 15316
rect 22764 15262 22766 15314
rect 22766 15262 22818 15314
rect 22818 15262 22820 15314
rect 22764 15260 22820 15262
rect 22988 16492 23044 16548
rect 24556 23378 24612 23380
rect 24556 23326 24558 23378
rect 24558 23326 24610 23378
rect 24610 23326 24612 23378
rect 24556 23324 24612 23326
rect 23548 20972 23604 21028
rect 23772 21196 23828 21252
rect 24332 22876 24388 22932
rect 23884 21084 23940 21140
rect 23772 20914 23828 20916
rect 23772 20862 23774 20914
rect 23774 20862 23826 20914
rect 23826 20862 23828 20914
rect 23772 20860 23828 20862
rect 24332 21586 24388 21588
rect 24332 21534 24334 21586
rect 24334 21534 24386 21586
rect 24386 21534 24388 21586
rect 24332 21532 24388 21534
rect 24444 22204 24500 22260
rect 24220 21474 24276 21476
rect 24220 21422 24222 21474
rect 24222 21422 24274 21474
rect 24274 21422 24276 21474
rect 24220 21420 24276 21422
rect 25340 24332 25396 24388
rect 25228 24220 25284 24276
rect 25004 23826 25060 23828
rect 25004 23774 25006 23826
rect 25006 23774 25058 23826
rect 25058 23774 25060 23826
rect 25004 23772 25060 23774
rect 24892 23660 24948 23716
rect 24780 22370 24836 22372
rect 24780 22318 24782 22370
rect 24782 22318 24834 22370
rect 24834 22318 24836 22370
rect 24780 22316 24836 22318
rect 24668 21868 24724 21924
rect 24556 21308 24612 21364
rect 24668 21586 24724 21588
rect 24668 21534 24670 21586
rect 24670 21534 24722 21586
rect 24722 21534 24724 21586
rect 24668 21532 24724 21534
rect 24108 20860 24164 20916
rect 23772 20188 23828 20244
rect 23660 20076 23716 20132
rect 23660 19404 23716 19460
rect 23660 18844 23716 18900
rect 23436 17554 23492 17556
rect 23436 17502 23438 17554
rect 23438 17502 23490 17554
rect 23490 17502 23492 17554
rect 23436 17500 23492 17502
rect 23660 17724 23716 17780
rect 23772 17666 23828 17668
rect 23772 17614 23774 17666
rect 23774 17614 23826 17666
rect 23826 17614 23828 17666
rect 23772 17612 23828 17614
rect 23212 16882 23268 16884
rect 23212 16830 23214 16882
rect 23214 16830 23266 16882
rect 23266 16830 23268 16882
rect 23212 16828 23268 16830
rect 23548 16716 23604 16772
rect 23212 16098 23268 16100
rect 23212 16046 23214 16098
rect 23214 16046 23266 16098
rect 23266 16046 23268 16098
rect 23212 16044 23268 16046
rect 23100 15932 23156 15988
rect 23100 15372 23156 15428
rect 22988 14530 23044 14532
rect 22988 14478 22990 14530
rect 22990 14478 23042 14530
rect 23042 14478 23044 14530
rect 22988 14476 23044 14478
rect 22652 13356 22708 13412
rect 22764 13244 22820 13300
rect 23436 15820 23492 15876
rect 23324 14476 23380 14532
rect 23436 14252 23492 14308
rect 23324 13356 23380 13412
rect 22652 12236 22708 12292
rect 22428 11340 22484 11396
rect 22540 12124 22596 12180
rect 22204 9212 22260 9268
rect 22092 9100 22148 9156
rect 21980 8428 22036 8484
rect 22092 8876 22148 8932
rect 21756 6188 21812 6244
rect 22204 8764 22260 8820
rect 22092 5964 22148 6020
rect 22316 8204 22372 8260
rect 22764 9884 22820 9940
rect 23436 12908 23492 12964
rect 23772 17276 23828 17332
rect 24108 20188 24164 20244
rect 25564 23826 25620 23828
rect 25564 23774 25566 23826
rect 25566 23774 25618 23826
rect 25618 23774 25620 23826
rect 25564 23772 25620 23774
rect 25340 23714 25396 23716
rect 25340 23662 25342 23714
rect 25342 23662 25394 23714
rect 25394 23662 25396 23714
rect 25340 23660 25396 23662
rect 25676 23324 25732 23380
rect 26460 23772 26516 23828
rect 26124 23324 26180 23380
rect 26124 23042 26180 23044
rect 26124 22990 26126 23042
rect 26126 22990 26178 23042
rect 26178 22990 26180 23042
rect 26124 22988 26180 22990
rect 25340 22930 25396 22932
rect 25340 22878 25342 22930
rect 25342 22878 25394 22930
rect 25394 22878 25396 22930
rect 25340 22876 25396 22878
rect 24892 20524 24948 20580
rect 23884 16770 23940 16772
rect 23884 16718 23886 16770
rect 23886 16718 23938 16770
rect 23938 16718 23940 16770
rect 23884 16716 23940 16718
rect 24108 19852 24164 19908
rect 24332 19740 24388 19796
rect 24780 19628 24836 19684
rect 24332 19458 24388 19460
rect 24332 19406 24334 19458
rect 24334 19406 24386 19458
rect 24386 19406 24388 19458
rect 24332 19404 24388 19406
rect 24332 18956 24388 19012
rect 24444 18674 24500 18676
rect 24444 18622 24446 18674
rect 24446 18622 24498 18674
rect 24498 18622 24500 18674
rect 24444 18620 24500 18622
rect 25452 22258 25508 22260
rect 25452 22206 25454 22258
rect 25454 22206 25506 22258
rect 25506 22206 25508 22258
rect 25452 22204 25508 22206
rect 25228 22146 25284 22148
rect 25228 22094 25230 22146
rect 25230 22094 25282 22146
rect 25282 22094 25284 22146
rect 25228 22092 25284 22094
rect 25116 21868 25172 21924
rect 25116 21196 25172 21252
rect 25116 19964 25172 20020
rect 25340 21810 25396 21812
rect 25340 21758 25342 21810
rect 25342 21758 25394 21810
rect 25394 21758 25396 21810
rect 25340 21756 25396 21758
rect 25340 21532 25396 21588
rect 26236 21644 26292 21700
rect 25788 21586 25844 21588
rect 25788 21534 25790 21586
rect 25790 21534 25842 21586
rect 25842 21534 25844 21586
rect 25788 21532 25844 21534
rect 26124 21420 26180 21476
rect 24108 17612 24164 17668
rect 24220 17500 24276 17556
rect 24108 16658 24164 16660
rect 24108 16606 24110 16658
rect 24110 16606 24162 16658
rect 24162 16606 24164 16658
rect 24108 16604 24164 16606
rect 24332 17836 24388 17892
rect 24780 17442 24836 17444
rect 24780 17390 24782 17442
rect 24782 17390 24834 17442
rect 24834 17390 24836 17442
rect 24780 17388 24836 17390
rect 23212 12066 23268 12068
rect 23212 12014 23214 12066
rect 23214 12014 23266 12066
rect 23266 12014 23268 12066
rect 23212 12012 23268 12014
rect 23324 12796 23380 12852
rect 22988 11340 23044 11396
rect 23100 9938 23156 9940
rect 23100 9886 23102 9938
rect 23102 9886 23154 9938
rect 23154 9886 23156 9938
rect 23100 9884 23156 9886
rect 22988 9660 23044 9716
rect 22764 9266 22820 9268
rect 22764 9214 22766 9266
rect 22766 9214 22818 9266
rect 22818 9214 22820 9266
rect 22764 9212 22820 9214
rect 22764 8764 22820 8820
rect 22540 7980 22596 8036
rect 23100 8258 23156 8260
rect 23100 8206 23102 8258
rect 23102 8206 23154 8258
rect 23154 8206 23156 8258
rect 23100 8204 23156 8206
rect 23772 13916 23828 13972
rect 23772 12796 23828 12852
rect 23884 12124 23940 12180
rect 23324 9154 23380 9156
rect 23324 9102 23326 9154
rect 23326 9102 23378 9154
rect 23378 9102 23380 9154
rect 23324 9100 23380 9102
rect 22540 6802 22596 6804
rect 22540 6750 22542 6802
rect 22542 6750 22594 6802
rect 22594 6750 22596 6802
rect 22540 6748 22596 6750
rect 22092 5628 22148 5684
rect 22540 5234 22596 5236
rect 22540 5182 22542 5234
rect 22542 5182 22594 5234
rect 22594 5182 22596 5234
rect 22540 5180 22596 5182
rect 21756 4172 21812 4228
rect 22428 4060 22484 4116
rect 22764 3612 22820 3668
rect 19068 3276 19124 3332
rect 22988 5964 23044 6020
rect 23100 5906 23156 5908
rect 23100 5854 23102 5906
rect 23102 5854 23154 5906
rect 23154 5854 23156 5906
rect 23100 5852 23156 5854
rect 23436 8764 23492 8820
rect 23436 7980 23492 8036
rect 23660 9042 23716 9044
rect 23660 8990 23662 9042
rect 23662 8990 23714 9042
rect 23714 8990 23716 9042
rect 23660 8988 23716 8990
rect 23884 11004 23940 11060
rect 23884 10556 23940 10612
rect 24108 13244 24164 13300
rect 24332 16380 24388 16436
rect 24780 17052 24836 17108
rect 24780 15932 24836 15988
rect 24332 15314 24388 15316
rect 24332 15262 24334 15314
rect 24334 15262 24386 15314
rect 24386 15262 24388 15314
rect 24332 15260 24388 15262
rect 24444 14364 24500 14420
rect 24668 14588 24724 14644
rect 25900 21196 25956 21252
rect 25676 20690 25732 20692
rect 25676 20638 25678 20690
rect 25678 20638 25730 20690
rect 25730 20638 25732 20690
rect 25676 20636 25732 20638
rect 25340 19516 25396 19572
rect 25340 19292 25396 19348
rect 25676 19740 25732 19796
rect 25788 19068 25844 19124
rect 25900 18844 25956 18900
rect 25788 18620 25844 18676
rect 26236 20524 26292 20580
rect 27468 26178 27524 26180
rect 27468 26126 27470 26178
rect 27470 26126 27522 26178
rect 27522 26126 27524 26178
rect 27468 26124 27524 26126
rect 26908 26012 26964 26068
rect 27244 26012 27300 26068
rect 28364 26066 28420 26068
rect 28364 26014 28366 26066
rect 28366 26014 28418 26066
rect 28418 26014 28420 26066
rect 28364 26012 28420 26014
rect 27916 25676 27972 25732
rect 30940 26348 30996 26404
rect 34300 30156 34356 30212
rect 33180 27692 33236 27748
rect 33628 29426 33684 29428
rect 33628 29374 33630 29426
rect 33630 29374 33682 29426
rect 33682 29374 33684 29426
rect 33628 29372 33684 29374
rect 36876 32674 36932 32676
rect 36876 32622 36878 32674
rect 36878 32622 36930 32674
rect 36930 32622 36932 32674
rect 36876 32620 36932 32622
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34748 30210 34804 30212
rect 34748 30158 34750 30210
rect 34750 30158 34802 30210
rect 34802 30158 34804 30210
rect 34748 30156 34804 30158
rect 35532 30210 35588 30212
rect 35532 30158 35534 30210
rect 35534 30158 35586 30210
rect 35586 30158 35588 30210
rect 35532 30156 35588 30158
rect 34860 30098 34916 30100
rect 34860 30046 34862 30098
rect 34862 30046 34914 30098
rect 34914 30046 34916 30098
rect 34860 30044 34916 30046
rect 36204 30322 36260 30324
rect 36204 30270 36206 30322
rect 36206 30270 36258 30322
rect 36258 30270 36260 30322
rect 36204 30268 36260 30270
rect 37324 33292 37380 33348
rect 38108 34354 38164 34356
rect 38108 34302 38110 34354
rect 38110 34302 38162 34354
rect 38162 34302 38164 34354
rect 38108 34300 38164 34302
rect 38556 37378 38612 37380
rect 38556 37326 38558 37378
rect 38558 37326 38610 37378
rect 38610 37326 38612 37378
rect 38556 37324 38612 37326
rect 39676 42140 39732 42196
rect 40236 42140 40292 42196
rect 39564 40962 39620 40964
rect 39564 40910 39566 40962
rect 39566 40910 39618 40962
rect 39618 40910 39620 40962
rect 39564 40908 39620 40910
rect 39116 39676 39172 39732
rect 39452 40514 39508 40516
rect 39452 40462 39454 40514
rect 39454 40462 39506 40514
rect 39506 40462 39508 40514
rect 39452 40460 39508 40462
rect 39900 41746 39956 41748
rect 39900 41694 39902 41746
rect 39902 41694 39954 41746
rect 39954 41694 39956 41746
rect 39900 41692 39956 41694
rect 39788 40460 39844 40516
rect 39564 40348 39620 40404
rect 39228 40124 39284 40180
rect 41244 44940 41300 44996
rect 41804 46674 41860 46676
rect 41804 46622 41806 46674
rect 41806 46622 41858 46674
rect 41858 46622 41860 46674
rect 41804 46620 41860 46622
rect 41356 44156 41412 44212
rect 41916 44156 41972 44212
rect 41020 44044 41076 44100
rect 41244 42364 41300 42420
rect 41020 41692 41076 41748
rect 40684 40012 40740 40068
rect 39564 39340 39620 39396
rect 40572 39340 40628 39396
rect 39788 39058 39844 39060
rect 39788 39006 39790 39058
rect 39790 39006 39842 39058
rect 39842 39006 39844 39058
rect 39788 39004 39844 39006
rect 39340 37378 39396 37380
rect 39340 37326 39342 37378
rect 39342 37326 39394 37378
rect 39394 37326 39396 37378
rect 39340 37324 39396 37326
rect 39788 37324 39844 37380
rect 39564 37266 39620 37268
rect 39564 37214 39566 37266
rect 39566 37214 39618 37266
rect 39618 37214 39620 37266
rect 39564 37212 39620 37214
rect 40012 37154 40068 37156
rect 40012 37102 40014 37154
rect 40014 37102 40066 37154
rect 40066 37102 40068 37154
rect 40012 37100 40068 37102
rect 39900 36988 39956 37044
rect 39116 36482 39172 36484
rect 39116 36430 39118 36482
rect 39118 36430 39170 36482
rect 39170 36430 39172 36482
rect 39116 36428 39172 36430
rect 40012 36652 40068 36708
rect 38892 36092 38948 36148
rect 38780 35868 38836 35924
rect 39676 35922 39732 35924
rect 39676 35870 39678 35922
rect 39678 35870 39730 35922
rect 39730 35870 39732 35922
rect 39676 35868 39732 35870
rect 40124 36428 40180 36484
rect 40012 34972 40068 35028
rect 41356 40460 41412 40516
rect 41580 40402 41636 40404
rect 41580 40350 41582 40402
rect 41582 40350 41634 40402
rect 41634 40350 41636 40402
rect 41580 40348 41636 40350
rect 41244 40012 41300 40068
rect 40796 39900 40852 39956
rect 43148 48300 43204 48356
rect 42588 46674 42644 46676
rect 42588 46622 42590 46674
rect 42590 46622 42642 46674
rect 42642 46622 42644 46674
rect 42588 46620 42644 46622
rect 46060 51436 46116 51492
rect 47180 53730 47236 53732
rect 47180 53678 47182 53730
rect 47182 53678 47234 53730
rect 47234 53678 47236 53730
rect 47180 53676 47236 53678
rect 49084 55020 49140 55076
rect 49308 54460 49364 54516
rect 47852 53676 47908 53732
rect 46844 51436 46900 51492
rect 45500 50876 45556 50932
rect 44492 50316 44548 50372
rect 45164 50428 45220 50484
rect 47404 51490 47460 51492
rect 47404 51438 47406 51490
rect 47406 51438 47458 51490
rect 47458 51438 47460 51490
rect 47404 51436 47460 51438
rect 46620 50428 46676 50484
rect 47068 50428 47124 50484
rect 45388 49586 45444 49588
rect 45388 49534 45390 49586
rect 45390 49534 45442 49586
rect 45442 49534 45444 49586
rect 45388 49532 45444 49534
rect 43596 49138 43652 49140
rect 43596 49086 43598 49138
rect 43598 49086 43650 49138
rect 43650 49086 43652 49138
rect 43596 49084 43652 49086
rect 46172 49532 46228 49588
rect 43932 48914 43988 48916
rect 43932 48862 43934 48914
rect 43934 48862 43986 48914
rect 43986 48862 43988 48914
rect 43932 48860 43988 48862
rect 43596 48748 43652 48804
rect 43484 47068 43540 47124
rect 42700 45330 42756 45332
rect 42700 45278 42702 45330
rect 42702 45278 42754 45330
rect 42754 45278 42756 45330
rect 42700 45276 42756 45278
rect 42252 45106 42308 45108
rect 42252 45054 42254 45106
rect 42254 45054 42306 45106
rect 42306 45054 42308 45106
rect 42252 45052 42308 45054
rect 42364 44994 42420 44996
rect 42364 44942 42366 44994
rect 42366 44942 42418 44994
rect 42418 44942 42420 44994
rect 42364 44940 42420 44942
rect 42028 42754 42084 42756
rect 42028 42702 42030 42754
rect 42030 42702 42082 42754
rect 42082 42702 42084 42754
rect 42028 42700 42084 42702
rect 44156 48802 44212 48804
rect 44156 48750 44158 48802
rect 44158 48750 44210 48802
rect 44210 48750 44212 48802
rect 44156 48748 44212 48750
rect 43932 48524 43988 48580
rect 44940 48466 44996 48468
rect 44940 48414 44942 48466
rect 44942 48414 44994 48466
rect 44994 48414 44996 48466
rect 44940 48412 44996 48414
rect 44044 48354 44100 48356
rect 44044 48302 44046 48354
rect 44046 48302 44098 48354
rect 44098 48302 44100 48354
rect 44044 48300 44100 48302
rect 44604 48300 44660 48356
rect 44156 46786 44212 46788
rect 44156 46734 44158 46786
rect 44158 46734 44210 46786
rect 44210 46734 44212 46786
rect 44156 46732 44212 46734
rect 43820 45890 43876 45892
rect 43820 45838 43822 45890
rect 43822 45838 43874 45890
rect 43874 45838 43876 45890
rect 43820 45836 43876 45838
rect 43708 45778 43764 45780
rect 43708 45726 43710 45778
rect 43710 45726 43762 45778
rect 43762 45726 43764 45778
rect 43708 45724 43764 45726
rect 42700 44210 42756 44212
rect 42700 44158 42702 44210
rect 42702 44158 42754 44210
rect 42754 44158 42756 44210
rect 42700 44156 42756 44158
rect 43148 43314 43204 43316
rect 43148 43262 43150 43314
rect 43150 43262 43202 43314
rect 43202 43262 43204 43314
rect 43148 43260 43204 43262
rect 43148 42866 43204 42868
rect 43148 42814 43150 42866
rect 43150 42814 43202 42866
rect 43202 42814 43204 42866
rect 43148 42812 43204 42814
rect 42140 42364 42196 42420
rect 43260 42364 43316 42420
rect 42476 41692 42532 41748
rect 41916 39900 41972 39956
rect 42028 40460 42084 40516
rect 41804 39564 41860 39620
rect 41468 39394 41524 39396
rect 41468 39342 41470 39394
rect 41470 39342 41522 39394
rect 41522 39342 41524 39394
rect 41468 39340 41524 39342
rect 41244 39058 41300 39060
rect 41244 39006 41246 39058
rect 41246 39006 41298 39058
rect 41298 39006 41300 39058
rect 41244 39004 41300 39006
rect 43148 40012 43204 40068
rect 42140 39618 42196 39620
rect 42140 39566 42142 39618
rect 42142 39566 42194 39618
rect 42194 39566 42196 39618
rect 42140 39564 42196 39566
rect 43484 40012 43540 40068
rect 42812 39340 42868 39396
rect 41580 38780 41636 38836
rect 42140 38610 42196 38612
rect 42140 38558 42142 38610
rect 42142 38558 42194 38610
rect 42194 38558 42196 38610
rect 42140 38556 42196 38558
rect 43484 39788 43540 39844
rect 43036 38946 43092 38948
rect 43036 38894 43038 38946
rect 43038 38894 43090 38946
rect 43090 38894 43092 38946
rect 43036 38892 43092 38894
rect 42476 37938 42532 37940
rect 42476 37886 42478 37938
rect 42478 37886 42530 37938
rect 42530 37886 42532 37938
rect 42476 37884 42532 37886
rect 41916 37490 41972 37492
rect 41916 37438 41918 37490
rect 41918 37438 41970 37490
rect 41970 37438 41972 37490
rect 41916 37436 41972 37438
rect 40908 37266 40964 37268
rect 40908 37214 40910 37266
rect 40910 37214 40962 37266
rect 40962 37214 40964 37266
rect 40908 37212 40964 37214
rect 41804 37100 41860 37156
rect 41132 36988 41188 37044
rect 42812 36876 42868 36932
rect 40908 36482 40964 36484
rect 40908 36430 40910 36482
rect 40910 36430 40962 36482
rect 40962 36430 40964 36482
rect 40908 36428 40964 36430
rect 41580 36370 41636 36372
rect 41580 36318 41582 36370
rect 41582 36318 41634 36370
rect 41634 36318 41636 36370
rect 41580 36316 41636 36318
rect 41916 35980 41972 36036
rect 42028 35868 42084 35924
rect 42812 36482 42868 36484
rect 42812 36430 42814 36482
rect 42814 36430 42866 36482
rect 42866 36430 42868 36482
rect 42812 36428 42868 36430
rect 40012 34802 40068 34804
rect 40012 34750 40014 34802
rect 40014 34750 40066 34802
rect 40066 34750 40068 34802
rect 40012 34748 40068 34750
rect 39116 34130 39172 34132
rect 39116 34078 39118 34130
rect 39118 34078 39170 34130
rect 39170 34078 39172 34130
rect 39116 34076 39172 34078
rect 39788 34130 39844 34132
rect 39788 34078 39790 34130
rect 39790 34078 39842 34130
rect 39842 34078 39844 34130
rect 39788 34076 39844 34078
rect 38220 33404 38276 33460
rect 38668 33964 38724 34020
rect 37212 32674 37268 32676
rect 37212 32622 37214 32674
rect 37214 32622 37266 32674
rect 37266 32622 37268 32674
rect 37212 32620 37268 32622
rect 38332 32674 38388 32676
rect 38332 32622 38334 32674
rect 38334 32622 38386 32674
rect 38386 32622 38388 32674
rect 38332 32620 38388 32622
rect 38220 32562 38276 32564
rect 38220 32510 38222 32562
rect 38222 32510 38274 32562
rect 38274 32510 38276 32562
rect 38220 32508 38276 32510
rect 37884 32396 37940 32452
rect 40348 34076 40404 34132
rect 41132 34130 41188 34132
rect 41132 34078 41134 34130
rect 41134 34078 41186 34130
rect 41186 34078 41188 34130
rect 41132 34076 41188 34078
rect 40908 33964 40964 34020
rect 40348 33234 40404 33236
rect 40348 33182 40350 33234
rect 40350 33182 40402 33234
rect 40402 33182 40404 33234
rect 40348 33180 40404 33182
rect 41356 33180 41412 33236
rect 43820 42476 43876 42532
rect 44940 48242 44996 48244
rect 44940 48190 44942 48242
rect 44942 48190 44994 48242
rect 44994 48190 44996 48242
rect 44940 48188 44996 48190
rect 44156 45500 44212 45556
rect 43820 40236 43876 40292
rect 43932 39618 43988 39620
rect 43932 39566 43934 39618
rect 43934 39566 43986 39618
rect 43986 39566 43988 39618
rect 43932 39564 43988 39566
rect 43820 39340 43876 39396
rect 44044 38892 44100 38948
rect 43596 38780 43652 38836
rect 43260 38722 43316 38724
rect 43260 38670 43262 38722
rect 43262 38670 43314 38722
rect 43314 38670 43316 38722
rect 43260 38668 43316 38670
rect 43932 38556 43988 38612
rect 43820 36540 43876 36596
rect 43036 36204 43092 36260
rect 43708 35980 43764 36036
rect 44044 36482 44100 36484
rect 44044 36430 44046 36482
rect 44046 36430 44098 36482
rect 44098 36430 44100 36482
rect 44044 36428 44100 36430
rect 45612 48188 45668 48244
rect 47964 50540 48020 50596
rect 46060 48802 46116 48804
rect 46060 48750 46062 48802
rect 46062 48750 46114 48802
rect 46114 48750 46116 48802
rect 46060 48748 46116 48750
rect 48636 50594 48692 50596
rect 48636 50542 48638 50594
rect 48638 50542 48690 50594
rect 48690 50542 48692 50594
rect 48636 50540 48692 50542
rect 49644 55410 49700 55412
rect 49644 55358 49646 55410
rect 49646 55358 49698 55410
rect 49698 55358 49700 55410
rect 49644 55356 49700 55358
rect 49980 55020 50036 55076
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 52220 56306 52276 56308
rect 52220 56254 52222 56306
rect 52222 56254 52274 56306
rect 52274 56254 52276 56306
rect 52220 56252 52276 56254
rect 51212 56082 51268 56084
rect 51212 56030 51214 56082
rect 51214 56030 51266 56082
rect 51266 56030 51268 56082
rect 51212 56028 51268 56030
rect 53116 56252 53172 56308
rect 54124 56306 54180 56308
rect 54124 56254 54126 56306
rect 54126 56254 54178 56306
rect 54178 56254 54180 56306
rect 54124 56252 54180 56254
rect 54460 56252 54516 56308
rect 55468 56306 55524 56308
rect 55468 56254 55470 56306
rect 55470 56254 55522 56306
rect 55522 56254 55524 56306
rect 55468 56252 55524 56254
rect 55132 55916 55188 55972
rect 55916 55970 55972 55972
rect 55916 55918 55918 55970
rect 55918 55918 55970 55970
rect 55970 55918 55972 55970
rect 55916 55916 55972 55918
rect 58156 55858 58212 55860
rect 58156 55806 58158 55858
rect 58158 55806 58210 55858
rect 58210 55806 58212 55858
rect 58156 55804 58212 55806
rect 52444 55356 52500 55412
rect 53676 55410 53732 55412
rect 53676 55358 53678 55410
rect 53678 55358 53730 55410
rect 53730 55358 53732 55410
rect 53676 55356 53732 55358
rect 51100 54796 51156 54852
rect 50092 54460 50148 54516
rect 52332 54796 52388 54852
rect 50876 54124 50932 54180
rect 50092 53730 50148 53732
rect 50092 53678 50094 53730
rect 50094 53678 50146 53730
rect 50146 53678 50148 53730
rect 50092 53676 50148 53678
rect 49644 53564 49700 53620
rect 50316 53506 50372 53508
rect 50316 53454 50318 53506
rect 50318 53454 50370 53506
rect 50370 53454 50372 53506
rect 50316 53452 50372 53454
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 49196 53004 49252 53060
rect 50652 53058 50708 53060
rect 50652 53006 50654 53058
rect 50654 53006 50706 53058
rect 50706 53006 50708 53058
rect 50652 53004 50708 53006
rect 50988 53730 51044 53732
rect 50988 53678 50990 53730
rect 50990 53678 51042 53730
rect 51042 53678 51044 53730
rect 50988 53676 51044 53678
rect 51660 53618 51716 53620
rect 51660 53566 51662 53618
rect 51662 53566 51714 53618
rect 51714 53566 51716 53618
rect 51660 53564 51716 53566
rect 52668 53618 52724 53620
rect 52668 53566 52670 53618
rect 52670 53566 52722 53618
rect 52722 53566 52724 53618
rect 52668 53564 52724 53566
rect 57708 55186 57764 55188
rect 57708 55134 57710 55186
rect 57710 55134 57762 55186
rect 57762 55134 57764 55186
rect 57708 55132 57764 55134
rect 58156 54460 58212 54516
rect 51324 53452 51380 53508
rect 51436 52162 51492 52164
rect 51436 52110 51438 52162
rect 51438 52110 51490 52162
rect 51490 52110 51492 52162
rect 51436 52108 51492 52110
rect 58156 52444 58212 52500
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50428 51212 50484 51268
rect 50652 50428 50708 50484
rect 51100 51996 51156 52052
rect 50988 50540 51044 50596
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49868 49810 49924 49812
rect 49868 49758 49870 49810
rect 49870 49758 49922 49810
rect 49922 49758 49924 49810
rect 49868 49756 49924 49758
rect 47740 49084 47796 49140
rect 47180 48748 47236 48804
rect 49084 48914 49140 48916
rect 49084 48862 49086 48914
rect 49086 48862 49138 48914
rect 49138 48862 49140 48914
rect 49084 48860 49140 48862
rect 47516 48748 47572 48804
rect 50092 49698 50148 49700
rect 50092 49646 50094 49698
rect 50094 49646 50146 49698
rect 50146 49646 50148 49698
rect 50092 49644 50148 49646
rect 51100 50482 51156 50484
rect 51100 50430 51102 50482
rect 51102 50430 51154 50482
rect 51154 50430 51156 50482
rect 51100 50428 51156 50430
rect 51212 51324 51268 51380
rect 50876 48914 50932 48916
rect 50876 48862 50878 48914
rect 50878 48862 50930 48914
rect 50930 48862 50932 48914
rect 50876 48860 50932 48862
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 49980 48412 50036 48468
rect 50988 48412 51044 48468
rect 45388 48018 45444 48020
rect 45388 47966 45390 48018
rect 45390 47966 45442 48018
rect 45442 47966 45444 48018
rect 45388 47964 45444 47966
rect 45500 47346 45556 47348
rect 45500 47294 45502 47346
rect 45502 47294 45554 47346
rect 45554 47294 45556 47346
rect 45500 47292 45556 47294
rect 45164 47068 45220 47124
rect 45052 46060 45108 46116
rect 45388 46674 45444 46676
rect 45388 46622 45390 46674
rect 45390 46622 45442 46674
rect 45442 46622 45444 46674
rect 45388 46620 45444 46622
rect 46396 47404 46452 47460
rect 49308 47570 49364 47572
rect 49308 47518 49310 47570
rect 49310 47518 49362 47570
rect 49362 47518 49364 47570
rect 49308 47516 49364 47518
rect 49532 47458 49588 47460
rect 49532 47406 49534 47458
rect 49534 47406 49586 47458
rect 49586 47406 49588 47458
rect 49532 47404 49588 47406
rect 50428 47404 50484 47460
rect 50652 47516 50708 47572
rect 46508 46786 46564 46788
rect 46508 46734 46510 46786
rect 46510 46734 46562 46786
rect 46562 46734 46564 46786
rect 46508 46732 46564 46734
rect 46732 46732 46788 46788
rect 46956 46620 47012 46676
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 51548 51212 51604 51268
rect 51660 50594 51716 50596
rect 51660 50542 51662 50594
rect 51662 50542 51714 50594
rect 51714 50542 51716 50594
rect 51660 50540 51716 50542
rect 52332 51324 52388 51380
rect 52892 50594 52948 50596
rect 52892 50542 52894 50594
rect 52894 50542 52946 50594
rect 52946 50542 52948 50594
rect 52892 50540 52948 50542
rect 57932 51100 57988 51156
rect 53900 50540 53956 50596
rect 55580 50594 55636 50596
rect 55580 50542 55582 50594
rect 55582 50542 55634 50594
rect 55634 50542 55636 50594
rect 55580 50540 55636 50542
rect 51884 50428 51940 50484
rect 52780 50482 52836 50484
rect 52780 50430 52782 50482
rect 52782 50430 52834 50482
rect 52834 50430 52836 50482
rect 52780 50428 52836 50430
rect 58156 50428 58212 50484
rect 58268 49084 58324 49140
rect 58156 48412 58212 48468
rect 53228 47404 53284 47460
rect 49868 46620 49924 46676
rect 50652 46674 50708 46676
rect 50652 46622 50654 46674
rect 50654 46622 50706 46674
rect 50706 46622 50708 46674
rect 50652 46620 50708 46622
rect 51324 46674 51380 46676
rect 51324 46622 51326 46674
rect 51326 46622 51378 46674
rect 51378 46622 51380 46674
rect 51324 46620 51380 46622
rect 48188 46562 48244 46564
rect 48188 46510 48190 46562
rect 48190 46510 48242 46562
rect 48242 46510 48244 46562
rect 48188 46508 48244 46510
rect 49532 46508 49588 46564
rect 46844 45890 46900 45892
rect 46844 45838 46846 45890
rect 46846 45838 46898 45890
rect 46898 45838 46900 45890
rect 46844 45836 46900 45838
rect 44940 45500 44996 45556
rect 44940 42812 44996 42868
rect 44828 42476 44884 42532
rect 44492 41746 44548 41748
rect 44492 41694 44494 41746
rect 44494 41694 44546 41746
rect 44546 41694 44548 41746
rect 44492 41692 44548 41694
rect 46172 44492 46228 44548
rect 45948 44322 46004 44324
rect 45948 44270 45950 44322
rect 45950 44270 46002 44322
rect 46002 44270 46004 44322
rect 45948 44268 46004 44270
rect 46396 44268 46452 44324
rect 46844 44322 46900 44324
rect 46844 44270 46846 44322
rect 46846 44270 46898 44322
rect 46898 44270 46900 44322
rect 46844 44268 46900 44270
rect 47404 44940 47460 44996
rect 50316 45890 50372 45892
rect 50316 45838 50318 45890
rect 50318 45838 50370 45890
rect 50370 45838 50372 45890
rect 50316 45836 50372 45838
rect 51660 46508 51716 46564
rect 51660 45890 51716 45892
rect 51660 45838 51662 45890
rect 51662 45838 51714 45890
rect 51714 45838 51716 45890
rect 51660 45836 51716 45838
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50092 44882 50148 44884
rect 50092 44830 50094 44882
rect 50094 44830 50146 44882
rect 50146 44830 50148 44882
rect 50092 44828 50148 44830
rect 47740 44716 47796 44772
rect 47516 44268 47572 44324
rect 49532 44716 49588 44772
rect 52444 45836 52500 45892
rect 53116 46562 53172 46564
rect 53116 46510 53118 46562
rect 53118 46510 53170 46562
rect 53170 46510 53172 46562
rect 53116 46508 53172 46510
rect 55580 47458 55636 47460
rect 55580 47406 55582 47458
rect 55582 47406 55634 47458
rect 55634 47406 55636 47458
rect 55580 47404 55636 47406
rect 57932 47068 57988 47124
rect 53340 46674 53396 46676
rect 53340 46622 53342 46674
rect 53342 46622 53394 46674
rect 53394 46622 53396 46674
rect 53340 46620 53396 46622
rect 50876 44828 50932 44884
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 53004 44268 53060 44324
rect 48300 43596 48356 43652
rect 49756 43650 49812 43652
rect 49756 43598 49758 43650
rect 49758 43598 49810 43650
rect 49810 43598 49812 43650
rect 49756 43596 49812 43598
rect 45052 42476 45108 42532
rect 45276 43314 45332 43316
rect 45276 43262 45278 43314
rect 45278 43262 45330 43314
rect 45330 43262 45332 43314
rect 45276 43260 45332 43262
rect 45276 42476 45332 42532
rect 45612 42530 45668 42532
rect 45612 42478 45614 42530
rect 45614 42478 45666 42530
rect 45666 42478 45668 42530
rect 45612 42476 45668 42478
rect 45836 41746 45892 41748
rect 45836 41694 45838 41746
rect 45838 41694 45890 41746
rect 45890 41694 45892 41746
rect 45836 41692 45892 41694
rect 46844 41916 46900 41972
rect 49868 43314 49924 43316
rect 49868 43262 49870 43314
rect 49870 43262 49922 43314
rect 49922 43262 49924 43314
rect 49868 43260 49924 43262
rect 47180 42194 47236 42196
rect 47180 42142 47182 42194
rect 47182 42142 47234 42194
rect 47234 42142 47236 42194
rect 47180 42140 47236 42142
rect 50092 42754 50148 42756
rect 50092 42702 50094 42754
rect 50094 42702 50146 42754
rect 50146 42702 50148 42754
rect 50092 42700 50148 42702
rect 49196 42140 49252 42196
rect 50652 43372 50708 43428
rect 48412 41916 48468 41972
rect 47404 41692 47460 41748
rect 45164 41244 45220 41300
rect 45948 41298 46004 41300
rect 45948 41246 45950 41298
rect 45950 41246 46002 41298
rect 46002 41246 46004 41298
rect 45948 41244 46004 41246
rect 51100 43484 51156 43540
rect 50764 42754 50820 42756
rect 50764 42702 50766 42754
rect 50766 42702 50818 42754
rect 50818 42702 50820 42754
rect 50764 42700 50820 42702
rect 50876 43260 50932 43316
rect 52332 43538 52388 43540
rect 52332 43486 52334 43538
rect 52334 43486 52386 43538
rect 52386 43486 52388 43538
rect 52332 43484 52388 43486
rect 52444 43426 52500 43428
rect 52444 43374 52446 43426
rect 52446 43374 52498 43426
rect 52498 43374 52500 43426
rect 52444 43372 52500 43374
rect 51212 43260 51268 43316
rect 55580 44322 55636 44324
rect 55580 44270 55582 44322
rect 55582 44270 55634 44322
rect 55634 44270 55636 44322
rect 55580 44268 55636 44270
rect 57932 43708 57988 43764
rect 51772 42700 51828 42756
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 55580 42754 55636 42756
rect 55580 42702 55582 42754
rect 55582 42702 55634 42754
rect 55634 42702 55636 42754
rect 55580 42700 55636 42702
rect 45052 40236 45108 40292
rect 48076 40908 48132 40964
rect 47852 40348 47908 40404
rect 45388 39618 45444 39620
rect 45388 39566 45390 39618
rect 45390 39566 45442 39618
rect 45442 39566 45444 39618
rect 45388 39564 45444 39566
rect 46284 39564 46340 39620
rect 45164 39506 45220 39508
rect 45164 39454 45166 39506
rect 45166 39454 45218 39506
rect 45218 39454 45220 39506
rect 45164 39452 45220 39454
rect 46620 39618 46676 39620
rect 46620 39566 46622 39618
rect 46622 39566 46674 39618
rect 46674 39566 46676 39618
rect 46620 39564 46676 39566
rect 46284 39058 46340 39060
rect 46284 39006 46286 39058
rect 46286 39006 46338 39058
rect 46338 39006 46340 39058
rect 46284 39004 46340 39006
rect 44268 38780 44324 38836
rect 46396 38834 46452 38836
rect 46396 38782 46398 38834
rect 46398 38782 46450 38834
rect 46450 38782 46452 38834
rect 46396 38780 46452 38782
rect 46508 38668 46564 38724
rect 46732 39004 46788 39060
rect 45836 37436 45892 37492
rect 47404 38834 47460 38836
rect 47404 38782 47406 38834
rect 47406 38782 47458 38834
rect 47458 38782 47460 38834
rect 47404 38780 47460 38782
rect 49084 40402 49140 40404
rect 49084 40350 49086 40402
rect 49086 40350 49138 40402
rect 49138 40350 49140 40402
rect 49084 40348 49140 40350
rect 57932 41692 57988 41748
rect 50428 41132 50484 41188
rect 49532 40908 49588 40964
rect 55580 41186 55636 41188
rect 55580 41134 55582 41186
rect 55582 41134 55634 41186
rect 55634 41134 55636 41186
rect 55580 41132 55636 41134
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 57932 40348 57988 40404
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 58268 39004 58324 39060
rect 46844 37436 46900 37492
rect 58156 38332 58212 38388
rect 49532 37996 49588 38052
rect 55580 38050 55636 38052
rect 55580 37998 55582 38050
rect 55582 37998 55634 38050
rect 55634 37998 55636 38050
rect 55580 37996 55636 37998
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 57932 37660 57988 37716
rect 50764 37604 50820 37606
rect 45612 36594 45668 36596
rect 45612 36542 45614 36594
rect 45614 36542 45666 36594
rect 45666 36542 45668 36594
rect 45612 36540 45668 36542
rect 47068 36594 47124 36596
rect 47068 36542 47070 36594
rect 47070 36542 47122 36594
rect 47122 36542 47124 36594
rect 47068 36540 47124 36542
rect 44156 36204 44212 36260
rect 44156 34972 44212 35028
rect 42140 33180 42196 33236
rect 38668 32732 38724 32788
rect 39004 32732 39060 32788
rect 39228 32562 39284 32564
rect 39228 32510 39230 32562
rect 39230 32510 39282 32562
rect 39282 32510 39284 32562
rect 39228 32508 39284 32510
rect 39676 32508 39732 32564
rect 38892 32396 38948 32452
rect 36988 30268 37044 30324
rect 35868 29708 35924 29764
rect 34412 29596 34468 29652
rect 34412 28588 34468 28644
rect 33404 27804 33460 27860
rect 31724 26348 31780 26404
rect 30828 26236 30884 26292
rect 29036 26178 29092 26180
rect 29036 26126 29038 26178
rect 29038 26126 29090 26178
rect 29090 26126 29092 26178
rect 29036 26124 29092 26126
rect 29708 25730 29764 25732
rect 29708 25678 29710 25730
rect 29710 25678 29762 25730
rect 29762 25678 29764 25730
rect 29708 25676 29764 25678
rect 30380 25676 30436 25732
rect 28252 25452 28308 25508
rect 29484 25506 29540 25508
rect 29484 25454 29486 25506
rect 29486 25454 29538 25506
rect 29538 25454 29540 25506
rect 29484 25452 29540 25454
rect 30716 25452 30772 25508
rect 27692 25282 27748 25284
rect 27692 25230 27694 25282
rect 27694 25230 27746 25282
rect 27746 25230 27748 25282
rect 27692 25228 27748 25230
rect 26684 23772 26740 23828
rect 27132 23938 27188 23940
rect 27132 23886 27134 23938
rect 27134 23886 27186 23938
rect 27186 23886 27188 23938
rect 27132 23884 27188 23886
rect 28028 24668 28084 24724
rect 27580 23826 27636 23828
rect 27580 23774 27582 23826
rect 27582 23774 27634 23826
rect 27634 23774 27636 23826
rect 27580 23772 27636 23774
rect 28700 25228 28756 25284
rect 28140 24220 28196 24276
rect 26908 23378 26964 23380
rect 26908 23326 26910 23378
rect 26910 23326 26962 23378
rect 26962 23326 26964 23378
rect 26908 23324 26964 23326
rect 27020 23154 27076 23156
rect 27020 23102 27022 23154
rect 27022 23102 27074 23154
rect 27074 23102 27076 23154
rect 27020 23100 27076 23102
rect 26684 22988 26740 23044
rect 27468 23212 27524 23268
rect 27692 23154 27748 23156
rect 27692 23102 27694 23154
rect 27694 23102 27746 23154
rect 27746 23102 27748 23154
rect 27692 23100 27748 23102
rect 28140 23324 28196 23380
rect 28028 22930 28084 22932
rect 28028 22878 28030 22930
rect 28030 22878 28082 22930
rect 28082 22878 28084 22930
rect 28028 22876 28084 22878
rect 26572 22316 26628 22372
rect 27804 22482 27860 22484
rect 27804 22430 27806 22482
rect 27806 22430 27858 22482
rect 27858 22430 27860 22482
rect 27804 22428 27860 22430
rect 26572 20748 26628 20804
rect 26572 20578 26628 20580
rect 26572 20526 26574 20578
rect 26574 20526 26626 20578
rect 26626 20526 26628 20578
rect 26572 20524 26628 20526
rect 26460 19234 26516 19236
rect 26460 19182 26462 19234
rect 26462 19182 26514 19234
rect 26514 19182 26516 19234
rect 26460 19180 26516 19182
rect 26348 18732 26404 18788
rect 25900 18508 25956 18564
rect 25564 18396 25620 18452
rect 25116 17666 25172 17668
rect 25116 17614 25118 17666
rect 25118 17614 25170 17666
rect 25170 17614 25172 17666
rect 25116 17612 25172 17614
rect 25228 17164 25284 17220
rect 25004 16492 25060 16548
rect 25676 16828 25732 16884
rect 25676 16380 25732 16436
rect 25340 16044 25396 16100
rect 24892 14418 24948 14420
rect 24892 14366 24894 14418
rect 24894 14366 24946 14418
rect 24946 14366 24948 14418
rect 24892 14364 24948 14366
rect 24668 13970 24724 13972
rect 24668 13918 24670 13970
rect 24670 13918 24722 13970
rect 24722 13918 24724 13970
rect 24668 13916 24724 13918
rect 24220 11340 24276 11396
rect 24108 10834 24164 10836
rect 24108 10782 24110 10834
rect 24110 10782 24162 10834
rect 24162 10782 24164 10834
rect 24108 10780 24164 10782
rect 24556 10780 24612 10836
rect 25788 16044 25844 16100
rect 25676 15596 25732 15652
rect 25228 13468 25284 13524
rect 25116 13356 25172 13412
rect 25004 13020 25060 13076
rect 25788 15148 25844 15204
rect 26236 17612 26292 17668
rect 26124 17052 26180 17108
rect 26684 19964 26740 20020
rect 26796 19404 26852 19460
rect 26684 19234 26740 19236
rect 26684 19182 26686 19234
rect 26686 19182 26738 19234
rect 26738 19182 26740 19234
rect 26684 19180 26740 19182
rect 27132 22258 27188 22260
rect 27132 22206 27134 22258
rect 27134 22206 27186 22258
rect 27186 22206 27188 22258
rect 27132 22204 27188 22206
rect 27132 21980 27188 22036
rect 27804 21868 27860 21924
rect 27692 21810 27748 21812
rect 27692 21758 27694 21810
rect 27694 21758 27746 21810
rect 27746 21758 27748 21810
rect 27692 21756 27748 21758
rect 27580 21308 27636 21364
rect 27244 20860 27300 20916
rect 27356 20578 27412 20580
rect 27356 20526 27358 20578
rect 27358 20526 27410 20578
rect 27410 20526 27412 20578
rect 27356 20524 27412 20526
rect 27132 19122 27188 19124
rect 27132 19070 27134 19122
rect 27134 19070 27186 19122
rect 27186 19070 27188 19122
rect 27132 19068 27188 19070
rect 26796 18396 26852 18452
rect 26908 18172 26964 18228
rect 26908 17388 26964 17444
rect 27244 17612 27300 17668
rect 27356 19516 27412 19572
rect 27692 19068 27748 19124
rect 30828 24722 30884 24724
rect 30828 24670 30830 24722
rect 30830 24670 30882 24722
rect 30882 24670 30884 24722
rect 30828 24668 30884 24670
rect 31500 25506 31556 25508
rect 31500 25454 31502 25506
rect 31502 25454 31554 25506
rect 31554 25454 31556 25506
rect 31500 25452 31556 25454
rect 32844 25506 32900 25508
rect 32844 25454 32846 25506
rect 32846 25454 32898 25506
rect 32898 25454 32900 25506
rect 32844 25452 32900 25454
rect 32060 25228 32116 25284
rect 31276 24668 31332 24724
rect 28364 23436 28420 23492
rect 30044 24108 30100 24164
rect 30268 23884 30324 23940
rect 30716 24108 30772 24164
rect 28476 23212 28532 23268
rect 28364 23154 28420 23156
rect 28364 23102 28366 23154
rect 28366 23102 28418 23154
rect 28418 23102 28420 23154
rect 28364 23100 28420 23102
rect 29484 23714 29540 23716
rect 29484 23662 29486 23714
rect 29486 23662 29538 23714
rect 29538 23662 29540 23714
rect 29484 23660 29540 23662
rect 28252 22652 28308 22708
rect 28364 22764 28420 22820
rect 28252 22370 28308 22372
rect 28252 22318 28254 22370
rect 28254 22318 28306 22370
rect 28306 22318 28308 22370
rect 28252 22316 28308 22318
rect 29148 22204 29204 22260
rect 27916 21084 27972 21140
rect 28028 20972 28084 21028
rect 27916 20412 27972 20468
rect 28364 20578 28420 20580
rect 28364 20526 28366 20578
rect 28366 20526 28418 20578
rect 28418 20526 28420 20578
rect 28364 20524 28420 20526
rect 29372 21532 29428 21588
rect 29372 21196 29428 21252
rect 28812 20412 28868 20468
rect 28140 19404 28196 19460
rect 28028 19010 28084 19012
rect 28028 18958 28030 19010
rect 28030 18958 28082 19010
rect 28082 18958 28084 19010
rect 28028 18956 28084 18958
rect 27692 18620 27748 18676
rect 28140 18732 28196 18788
rect 27580 18450 27636 18452
rect 27580 18398 27582 18450
rect 27582 18398 27634 18450
rect 27634 18398 27636 18450
rect 27580 18396 27636 18398
rect 27356 17388 27412 17444
rect 26460 16716 26516 16772
rect 26908 16268 26964 16324
rect 26572 16210 26628 16212
rect 26572 16158 26574 16210
rect 26574 16158 26626 16210
rect 26626 16158 26628 16210
rect 26572 16156 26628 16158
rect 26460 15932 26516 15988
rect 26684 16044 26740 16100
rect 26460 15596 26516 15652
rect 26124 15260 26180 15316
rect 25676 14476 25732 14532
rect 25452 13858 25508 13860
rect 25452 13806 25454 13858
rect 25454 13806 25506 13858
rect 25506 13806 25508 13858
rect 25452 13804 25508 13806
rect 25788 13804 25844 13860
rect 26012 14306 26068 14308
rect 26012 14254 26014 14306
rect 26014 14254 26066 14306
rect 26066 14254 26068 14306
rect 26012 14252 26068 14254
rect 25564 13244 25620 13300
rect 25452 12796 25508 12852
rect 25004 11788 25060 11844
rect 25116 11618 25172 11620
rect 25116 11566 25118 11618
rect 25118 11566 25170 11618
rect 25170 11566 25172 11618
rect 25116 11564 25172 11566
rect 24108 9436 24164 9492
rect 24220 9826 24276 9828
rect 24220 9774 24222 9826
rect 24222 9774 24274 9826
rect 24274 9774 24276 9826
rect 24220 9772 24276 9774
rect 24220 9100 24276 9156
rect 23884 8988 23940 9044
rect 23660 8652 23716 8708
rect 24108 7532 24164 7588
rect 24108 6524 24164 6580
rect 24220 7308 24276 7364
rect 23436 6188 23492 6244
rect 25004 10668 25060 10724
rect 24668 10444 24724 10500
rect 24892 10556 24948 10612
rect 24668 10220 24724 10276
rect 24780 10332 24836 10388
rect 24444 10108 24500 10164
rect 24668 9996 24724 10052
rect 24332 8204 24388 8260
rect 24556 8316 24612 8372
rect 24444 7474 24500 7476
rect 24444 7422 24446 7474
rect 24446 7422 24498 7474
rect 24498 7422 24500 7474
rect 24444 7420 24500 7422
rect 24444 6860 24500 6916
rect 24556 6076 24612 6132
rect 24332 5516 24388 5572
rect 24220 4620 24276 4676
rect 24332 5180 24388 5236
rect 23436 4060 23492 4116
rect 23996 4284 24052 4340
rect 23548 3554 23604 3556
rect 23548 3502 23550 3554
rect 23550 3502 23602 3554
rect 23602 3502 23604 3554
rect 23548 3500 23604 3502
rect 24444 4956 24500 5012
rect 23212 3442 23268 3444
rect 23212 3390 23214 3442
rect 23214 3390 23266 3442
rect 23266 3390 23268 3442
rect 23212 3388 23268 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22988 3276 23044 3332
rect 20412 3052 20468 3108
rect 19516 2940 19572 2996
rect 18956 2716 19012 2772
rect 25676 11900 25732 11956
rect 25564 10668 25620 10724
rect 25116 9826 25172 9828
rect 25116 9774 25118 9826
rect 25118 9774 25170 9826
rect 25170 9774 25172 9826
rect 25116 9772 25172 9774
rect 25564 10444 25620 10500
rect 25452 9884 25508 9940
rect 25228 8876 25284 8932
rect 25340 9548 25396 9604
rect 25340 8540 25396 8596
rect 25452 8764 25508 8820
rect 25228 8316 25284 8372
rect 25228 8092 25284 8148
rect 25340 7586 25396 7588
rect 25340 7534 25342 7586
rect 25342 7534 25394 7586
rect 25394 7534 25396 7586
rect 25340 7532 25396 7534
rect 25340 7250 25396 7252
rect 25340 7198 25342 7250
rect 25342 7198 25394 7250
rect 25394 7198 25396 7250
rect 25340 7196 25396 7198
rect 25228 6018 25284 6020
rect 25228 5966 25230 6018
rect 25230 5966 25282 6018
rect 25282 5966 25284 6018
rect 25228 5964 25284 5966
rect 26124 13244 26180 13300
rect 25900 11228 25956 11284
rect 26124 11676 26180 11732
rect 26124 11394 26180 11396
rect 26124 11342 26126 11394
rect 26126 11342 26178 11394
rect 26178 11342 26180 11394
rect 26124 11340 26180 11342
rect 26236 10332 26292 10388
rect 26572 15036 26628 15092
rect 26908 12962 26964 12964
rect 26908 12910 26910 12962
rect 26910 12910 26962 12962
rect 26962 12910 26964 12962
rect 26908 12908 26964 12910
rect 27132 16828 27188 16884
rect 28140 18284 28196 18340
rect 28364 18562 28420 18564
rect 28364 18510 28366 18562
rect 28366 18510 28418 18562
rect 28418 18510 28420 18562
rect 28364 18508 28420 18510
rect 27692 17388 27748 17444
rect 28140 17388 28196 17444
rect 28252 17724 28308 17780
rect 27580 16716 27636 16772
rect 27356 16492 27412 16548
rect 27468 16098 27524 16100
rect 27468 16046 27470 16098
rect 27470 16046 27522 16098
rect 27522 16046 27524 16098
rect 27468 16044 27524 16046
rect 27580 16268 27636 16324
rect 27356 15484 27412 15540
rect 27804 16882 27860 16884
rect 27804 16830 27806 16882
rect 27806 16830 27858 16882
rect 27858 16830 27860 16882
rect 27804 16828 27860 16830
rect 28140 15820 28196 15876
rect 27692 15314 27748 15316
rect 27692 15262 27694 15314
rect 27694 15262 27746 15314
rect 27746 15262 27748 15314
rect 27692 15260 27748 15262
rect 27356 14588 27412 14644
rect 27132 14418 27188 14420
rect 27132 14366 27134 14418
rect 27134 14366 27186 14418
rect 27186 14366 27188 14418
rect 27132 14364 27188 14366
rect 27468 14530 27524 14532
rect 27468 14478 27470 14530
rect 27470 14478 27522 14530
rect 27522 14478 27524 14530
rect 27468 14476 27524 14478
rect 27580 14924 27636 14980
rect 27356 13692 27412 13748
rect 27804 15036 27860 15092
rect 27692 14418 27748 14420
rect 27692 14366 27694 14418
rect 27694 14366 27746 14418
rect 27746 14366 27748 14418
rect 27692 14364 27748 14366
rect 27692 14028 27748 14084
rect 27916 14140 27972 14196
rect 28028 13916 28084 13972
rect 27132 12684 27188 12740
rect 26684 10610 26740 10612
rect 26684 10558 26686 10610
rect 26686 10558 26738 10610
rect 26738 10558 26740 10610
rect 26684 10556 26740 10558
rect 25676 8876 25732 8932
rect 25788 8258 25844 8260
rect 25788 8206 25790 8258
rect 25790 8206 25842 8258
rect 25842 8206 25844 8258
rect 25788 8204 25844 8206
rect 25788 7644 25844 7700
rect 25564 4172 25620 4228
rect 25788 5964 25844 6020
rect 26012 5628 26068 5684
rect 26684 9100 26740 9156
rect 26460 8876 26516 8932
rect 26236 8540 26292 8596
rect 26348 8146 26404 8148
rect 26348 8094 26350 8146
rect 26350 8094 26402 8146
rect 26402 8094 26404 8146
rect 26348 8092 26404 8094
rect 27020 11282 27076 11284
rect 27020 11230 27022 11282
rect 27022 11230 27074 11282
rect 27074 11230 27076 11282
rect 27020 11228 27076 11230
rect 27244 11228 27300 11284
rect 27244 9996 27300 10052
rect 27356 9884 27412 9940
rect 27020 9826 27076 9828
rect 27020 9774 27022 9826
rect 27022 9774 27074 9826
rect 27074 9774 27076 9826
rect 27020 9772 27076 9774
rect 27132 9042 27188 9044
rect 27132 8990 27134 9042
rect 27134 8990 27186 9042
rect 27186 8990 27188 9042
rect 27132 8988 27188 8990
rect 26908 8428 26964 8484
rect 26124 4844 26180 4900
rect 26460 5740 26516 5796
rect 26572 6972 26628 7028
rect 27020 7980 27076 8036
rect 26684 6748 26740 6804
rect 26684 6466 26740 6468
rect 26684 6414 26686 6466
rect 26686 6414 26738 6466
rect 26738 6414 26740 6466
rect 26684 6412 26740 6414
rect 26908 6412 26964 6468
rect 26796 6130 26852 6132
rect 26796 6078 26798 6130
rect 26798 6078 26850 6130
rect 26850 6078 26852 6130
rect 26796 6076 26852 6078
rect 28252 15426 28308 15428
rect 28252 15374 28254 15426
rect 28254 15374 28306 15426
rect 28306 15374 28308 15426
rect 28252 15372 28308 15374
rect 29372 20412 29428 20468
rect 28924 19516 28980 19572
rect 29036 18620 29092 18676
rect 28924 18508 28980 18564
rect 28588 15708 28644 15764
rect 28588 15372 28644 15428
rect 29036 18172 29092 18228
rect 30268 23660 30324 23716
rect 30604 23714 30660 23716
rect 30604 23662 30606 23714
rect 30606 23662 30658 23714
rect 30658 23662 30660 23714
rect 30604 23660 30660 23662
rect 30380 22988 30436 23044
rect 30268 22876 30324 22932
rect 29932 22316 29988 22372
rect 30044 22204 30100 22260
rect 29708 22092 29764 22148
rect 30156 20972 30212 21028
rect 30268 21420 30324 21476
rect 29596 20860 29652 20916
rect 29932 20578 29988 20580
rect 29932 20526 29934 20578
rect 29934 20526 29986 20578
rect 29986 20526 29988 20578
rect 29932 20524 29988 20526
rect 31164 23884 31220 23940
rect 31948 25004 32004 25060
rect 31724 23548 31780 23604
rect 31836 23212 31892 23268
rect 31052 22876 31108 22932
rect 31500 23154 31556 23156
rect 31500 23102 31502 23154
rect 31502 23102 31554 23154
rect 31554 23102 31556 23154
rect 31500 23100 31556 23102
rect 31388 22652 31444 22708
rect 31276 22594 31332 22596
rect 31276 22542 31278 22594
rect 31278 22542 31330 22594
rect 31330 22542 31332 22594
rect 31276 22540 31332 22542
rect 30940 22204 30996 22260
rect 30716 21980 30772 22036
rect 30828 21586 30884 21588
rect 30828 21534 30830 21586
rect 30830 21534 30882 21586
rect 30882 21534 30884 21586
rect 30828 21532 30884 21534
rect 31388 21644 31444 21700
rect 31052 21420 31108 21476
rect 31276 21362 31332 21364
rect 31276 21310 31278 21362
rect 31278 21310 31330 21362
rect 31330 21310 31332 21362
rect 31276 21308 31332 21310
rect 30380 20524 30436 20580
rect 30828 20972 30884 21028
rect 30268 20188 30324 20244
rect 30492 20300 30548 20356
rect 30156 19740 30212 19796
rect 29484 19234 29540 19236
rect 29484 19182 29486 19234
rect 29486 19182 29538 19234
rect 29538 19182 29540 19234
rect 29484 19180 29540 19182
rect 29596 18674 29652 18676
rect 29596 18622 29598 18674
rect 29598 18622 29650 18674
rect 29650 18622 29652 18674
rect 29596 18620 29652 18622
rect 28924 16268 28980 16324
rect 29036 17388 29092 17444
rect 28812 15932 28868 15988
rect 28700 15260 28756 15316
rect 29148 16940 29204 16996
rect 29148 16492 29204 16548
rect 29596 17164 29652 17220
rect 29372 17052 29428 17108
rect 29932 17052 29988 17108
rect 29484 16268 29540 16324
rect 28588 14924 28644 14980
rect 28252 14476 28308 14532
rect 28476 14476 28532 14532
rect 28476 13468 28532 13524
rect 28252 13244 28308 13300
rect 28252 13020 28308 13076
rect 28924 14140 28980 14196
rect 28028 12684 28084 12740
rect 27580 11452 27636 11508
rect 27804 12460 27860 12516
rect 27580 10834 27636 10836
rect 27580 10782 27582 10834
rect 27582 10782 27634 10834
rect 27634 10782 27636 10834
rect 27580 10780 27636 10782
rect 28252 12012 28308 12068
rect 28364 11954 28420 11956
rect 28364 11902 28366 11954
rect 28366 11902 28418 11954
rect 28418 11902 28420 11954
rect 28364 11900 28420 11902
rect 28588 11676 28644 11732
rect 28700 11564 28756 11620
rect 27916 9996 27972 10052
rect 28140 10498 28196 10500
rect 28140 10446 28142 10498
rect 28142 10446 28194 10498
rect 28194 10446 28196 10498
rect 28140 10444 28196 10446
rect 28700 11228 28756 11284
rect 28364 10780 28420 10836
rect 27356 6972 27412 7028
rect 27692 9266 27748 9268
rect 27692 9214 27694 9266
rect 27694 9214 27746 9266
rect 27746 9214 27748 9266
rect 27692 9212 27748 9214
rect 27692 7756 27748 7812
rect 28252 9826 28308 9828
rect 28252 9774 28254 9826
rect 28254 9774 28306 9826
rect 28306 9774 28308 9826
rect 28252 9772 28308 9774
rect 28028 9154 28084 9156
rect 28028 9102 28030 9154
rect 28030 9102 28082 9154
rect 28082 9102 28084 9154
rect 28028 9100 28084 9102
rect 28028 8258 28084 8260
rect 28028 8206 28030 8258
rect 28030 8206 28082 8258
rect 28082 8206 28084 8258
rect 28028 8204 28084 8206
rect 28028 7868 28084 7924
rect 27916 7644 27972 7700
rect 28140 7644 28196 7700
rect 28028 7532 28084 7588
rect 27916 7420 27972 7476
rect 27020 5964 27076 6020
rect 27244 6748 27300 6804
rect 27692 6860 27748 6916
rect 27244 6466 27300 6468
rect 27244 6414 27246 6466
rect 27246 6414 27298 6466
rect 27298 6414 27300 6466
rect 27244 6412 27300 6414
rect 27356 5852 27412 5908
rect 27468 6412 27524 6468
rect 26236 5516 26292 5572
rect 26348 5292 26404 5348
rect 26572 5234 26628 5236
rect 26572 5182 26574 5234
rect 26574 5182 26626 5234
rect 26626 5182 26628 5234
rect 26572 5180 26628 5182
rect 26572 4956 26628 5012
rect 26348 4844 26404 4900
rect 26236 4508 26292 4564
rect 26684 4284 26740 4340
rect 24668 2268 24724 2324
rect 18844 1596 18900 1652
rect 27356 5234 27412 5236
rect 27356 5182 27358 5234
rect 27358 5182 27410 5234
rect 27410 5182 27412 5234
rect 27356 5180 27412 5182
rect 27356 4844 27412 4900
rect 27244 4562 27300 4564
rect 27244 4510 27246 4562
rect 27246 4510 27298 4562
rect 27298 4510 27300 4562
rect 27244 4508 27300 4510
rect 27916 7084 27972 7140
rect 27804 6524 27860 6580
rect 27580 6018 27636 6020
rect 27580 5966 27582 6018
rect 27582 5966 27634 6018
rect 27634 5966 27636 6018
rect 27580 5964 27636 5966
rect 27804 5852 27860 5908
rect 27692 5628 27748 5684
rect 27468 4508 27524 4564
rect 28140 7420 28196 7476
rect 28140 7196 28196 7252
rect 28700 9772 28756 9828
rect 28924 10444 28980 10500
rect 28812 9212 28868 9268
rect 29148 14306 29204 14308
rect 29148 14254 29150 14306
rect 29150 14254 29202 14306
rect 29202 14254 29204 14306
rect 29148 14252 29204 14254
rect 29372 14028 29428 14084
rect 29148 10892 29204 10948
rect 28364 8316 28420 8372
rect 28252 5516 28308 5572
rect 29148 9100 29204 9156
rect 28588 7532 28644 7588
rect 28476 7196 28532 7252
rect 28476 5740 28532 5796
rect 27356 3666 27412 3668
rect 27356 3614 27358 3666
rect 27358 3614 27410 3666
rect 27410 3614 27412 3666
rect 27356 3612 27412 3614
rect 27804 3554 27860 3556
rect 27804 3502 27806 3554
rect 27806 3502 27858 3554
rect 27858 3502 27860 3554
rect 27804 3500 27860 3502
rect 28588 4732 28644 4788
rect 28812 6524 28868 6580
rect 29036 8092 29092 8148
rect 30380 19458 30436 19460
rect 30380 19406 30382 19458
rect 30382 19406 30434 19458
rect 30434 19406 30436 19458
rect 30380 19404 30436 19406
rect 30604 19628 30660 19684
rect 30268 18956 30324 19012
rect 30380 17836 30436 17892
rect 30492 18396 30548 18452
rect 30156 16940 30212 16996
rect 30268 17164 30324 17220
rect 29932 15708 29988 15764
rect 30156 15426 30212 15428
rect 30156 15374 30158 15426
rect 30158 15374 30210 15426
rect 30210 15374 30212 15426
rect 30156 15372 30212 15374
rect 29820 14588 29876 14644
rect 29708 14364 29764 14420
rect 29820 12178 29876 12180
rect 29820 12126 29822 12178
rect 29822 12126 29874 12178
rect 29874 12126 29876 12178
rect 29820 12124 29876 12126
rect 29708 12066 29764 12068
rect 29708 12014 29710 12066
rect 29710 12014 29762 12066
rect 29762 12014 29764 12066
rect 29708 12012 29764 12014
rect 29820 11676 29876 11732
rect 29372 10556 29428 10612
rect 29820 10220 29876 10276
rect 29372 8258 29428 8260
rect 29372 8206 29374 8258
rect 29374 8206 29426 8258
rect 29426 8206 29428 8258
rect 29372 8204 29428 8206
rect 29148 7474 29204 7476
rect 29148 7422 29150 7474
rect 29150 7422 29202 7474
rect 29202 7422 29204 7474
rect 29148 7420 29204 7422
rect 29148 5852 29204 5908
rect 28924 4732 28980 4788
rect 29036 5068 29092 5124
rect 28700 4172 28756 4228
rect 29260 4956 29316 5012
rect 29148 4284 29204 4340
rect 29484 4172 29540 4228
rect 29708 8428 29764 8484
rect 30156 14924 30212 14980
rect 31164 20636 31220 20692
rect 31724 21084 31780 21140
rect 31388 20524 31444 20580
rect 31164 20188 31220 20244
rect 32060 24722 32116 24724
rect 32060 24670 32062 24722
rect 32062 24670 32114 24722
rect 32114 24670 32116 24722
rect 32060 24668 32116 24670
rect 32620 24556 32676 24612
rect 32508 23266 32564 23268
rect 32508 23214 32510 23266
rect 32510 23214 32562 23266
rect 32562 23214 32564 23266
rect 32508 23212 32564 23214
rect 32172 23042 32228 23044
rect 32172 22990 32174 23042
rect 32174 22990 32226 23042
rect 32226 22990 32228 23042
rect 32172 22988 32228 22990
rect 32508 22652 32564 22708
rect 32284 21084 32340 21140
rect 31836 20412 31892 20468
rect 30716 17666 30772 17668
rect 30716 17614 30718 17666
rect 30718 17614 30770 17666
rect 30770 17614 30772 17666
rect 30716 17612 30772 17614
rect 30940 19906 30996 19908
rect 30940 19854 30942 19906
rect 30942 19854 30994 19906
rect 30994 19854 30996 19906
rect 30940 19852 30996 19854
rect 30940 18060 30996 18116
rect 31052 17836 31108 17892
rect 30492 17052 30548 17108
rect 30940 17500 30996 17556
rect 30380 15484 30436 15540
rect 30044 8316 30100 8372
rect 30268 13020 30324 13076
rect 29932 8258 29988 8260
rect 29932 8206 29934 8258
rect 29934 8206 29986 8258
rect 29986 8206 29988 8258
rect 29932 8204 29988 8206
rect 30828 16940 30884 16996
rect 31052 17052 31108 17108
rect 31836 20076 31892 20132
rect 31500 19234 31556 19236
rect 31500 19182 31502 19234
rect 31502 19182 31554 19234
rect 31554 19182 31556 19234
rect 31500 19180 31556 19182
rect 31724 17612 31780 17668
rect 31500 16828 31556 16884
rect 31164 15708 31220 15764
rect 31052 13746 31108 13748
rect 31052 13694 31054 13746
rect 31054 13694 31106 13746
rect 31106 13694 31108 13746
rect 31052 13692 31108 13694
rect 30716 12908 30772 12964
rect 30828 13580 30884 13636
rect 31052 13468 31108 13524
rect 30268 10610 30324 10612
rect 30268 10558 30270 10610
rect 30270 10558 30322 10610
rect 30322 10558 30324 10610
rect 30268 10556 30324 10558
rect 30492 11282 30548 11284
rect 30492 11230 30494 11282
rect 30494 11230 30546 11282
rect 30546 11230 30548 11282
rect 30492 11228 30548 11230
rect 30716 11228 30772 11284
rect 31052 10668 31108 10724
rect 30828 10444 30884 10500
rect 30604 8316 30660 8372
rect 30380 8034 30436 8036
rect 30380 7982 30382 8034
rect 30382 7982 30434 8034
rect 30434 7982 30436 8034
rect 30380 7980 30436 7982
rect 30604 8146 30660 8148
rect 30604 8094 30606 8146
rect 30606 8094 30658 8146
rect 30658 8094 30660 8146
rect 30604 8092 30660 8094
rect 30156 7532 30212 7588
rect 29708 5964 29764 6020
rect 30380 7474 30436 7476
rect 30380 7422 30382 7474
rect 30382 7422 30434 7474
rect 30434 7422 30436 7474
rect 30380 7420 30436 7422
rect 29932 5292 29988 5348
rect 29708 5068 29764 5124
rect 30044 5010 30100 5012
rect 30044 4958 30046 5010
rect 30046 4958 30098 5010
rect 30098 4958 30100 5010
rect 30044 4956 30100 4958
rect 30940 8988 30996 9044
rect 30940 7980 30996 8036
rect 30716 7644 30772 7700
rect 30716 7420 30772 7476
rect 31276 14700 31332 14756
rect 31388 14588 31444 14644
rect 31276 14530 31332 14532
rect 31276 14478 31278 14530
rect 31278 14478 31330 14530
rect 31330 14478 31332 14530
rect 31276 14476 31332 14478
rect 31388 12962 31444 12964
rect 31388 12910 31390 12962
rect 31390 12910 31442 12962
rect 31442 12910 31444 12962
rect 31388 12908 31444 12910
rect 31388 12738 31444 12740
rect 31388 12686 31390 12738
rect 31390 12686 31442 12738
rect 31442 12686 31444 12738
rect 31388 12684 31444 12686
rect 31388 12236 31444 12292
rect 31388 10892 31444 10948
rect 31612 14140 31668 14196
rect 32396 20018 32452 20020
rect 32396 19966 32398 20018
rect 32398 19966 32450 20018
rect 32450 19966 32452 20018
rect 32396 19964 32452 19966
rect 32172 19852 32228 19908
rect 32060 19404 32116 19460
rect 32956 24050 33012 24052
rect 32956 23998 32958 24050
rect 32958 23998 33010 24050
rect 33010 23998 33012 24050
rect 32956 23996 33012 23998
rect 33068 21698 33124 21700
rect 33068 21646 33070 21698
rect 33070 21646 33122 21698
rect 33122 21646 33124 21698
rect 33068 21644 33124 21646
rect 32844 20860 32900 20916
rect 33516 27692 33572 27748
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34972 27804 35028 27860
rect 36876 29708 36932 29764
rect 36988 28642 37044 28644
rect 36988 28590 36990 28642
rect 36990 28590 37042 28642
rect 37042 28590 37044 28642
rect 36988 28588 37044 28590
rect 38108 29708 38164 29764
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 38892 29426 38948 29428
rect 38892 29374 38894 29426
rect 38894 29374 38946 29426
rect 38946 29374 38948 29426
rect 38892 29372 38948 29374
rect 45836 36316 45892 36372
rect 46844 36316 46900 36372
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 46732 35810 46788 35812
rect 46732 35758 46734 35810
rect 46734 35758 46786 35810
rect 46786 35758 46788 35810
rect 46732 35756 46788 35758
rect 55580 35756 55636 35812
rect 57820 36316 57876 36372
rect 57932 35644 57988 35700
rect 45388 34860 45444 34916
rect 55580 34914 55636 34916
rect 55580 34862 55582 34914
rect 55582 34862 55634 34914
rect 55634 34862 55636 34914
rect 55580 34860 55636 34862
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 44156 34130 44212 34132
rect 44156 34078 44158 34130
rect 44158 34078 44210 34130
rect 44210 34078 44212 34130
rect 44156 34076 44212 34078
rect 43484 33964 43540 34020
rect 45388 34076 45444 34132
rect 44604 33964 44660 34020
rect 45276 33964 45332 34020
rect 45052 33346 45108 33348
rect 45052 33294 45054 33346
rect 45054 33294 45106 33346
rect 45106 33294 45108 33346
rect 45052 33292 45108 33294
rect 41916 31052 41972 31108
rect 58156 33628 58212 33684
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 58156 32956 58212 33012
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 57820 31106 57876 31108
rect 57820 31054 57822 31106
rect 57822 31054 57874 31106
rect 57874 31054 57876 31106
rect 57820 31052 57876 31054
rect 58156 30268 58212 30324
rect 41916 30044 41972 30100
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 41580 29426 41636 29428
rect 41580 29374 41582 29426
rect 41582 29374 41634 29426
rect 41634 29374 41636 29426
rect 41580 29372 41636 29374
rect 37996 27804 38052 27860
rect 37212 27020 37268 27076
rect 37772 27244 37828 27300
rect 34188 26012 34244 26068
rect 33852 25676 33908 25732
rect 33740 25228 33796 25284
rect 33628 24834 33684 24836
rect 33628 24782 33630 24834
rect 33630 24782 33682 24834
rect 33682 24782 33684 24834
rect 33628 24780 33684 24782
rect 33292 24722 33348 24724
rect 33292 24670 33294 24722
rect 33294 24670 33346 24722
rect 33346 24670 33348 24722
rect 33292 24668 33348 24670
rect 33292 23772 33348 23828
rect 33740 23042 33796 23044
rect 33740 22990 33742 23042
rect 33742 22990 33794 23042
rect 33794 22990 33796 23042
rect 33740 22988 33796 22990
rect 34076 25564 34132 25620
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34636 25676 34692 25732
rect 34300 24668 34356 24724
rect 33628 22428 33684 22484
rect 33964 23772 34020 23828
rect 33404 21810 33460 21812
rect 33404 21758 33406 21810
rect 33406 21758 33458 21810
rect 33458 21758 33460 21810
rect 33404 21756 33460 21758
rect 33292 20300 33348 20356
rect 32172 18284 32228 18340
rect 32172 18060 32228 18116
rect 31948 17724 32004 17780
rect 31836 17500 31892 17556
rect 32060 17164 32116 17220
rect 33180 18620 33236 18676
rect 33740 21644 33796 21700
rect 35532 25676 35588 25732
rect 35196 24780 35252 24836
rect 34860 24444 34916 24500
rect 34748 23772 34804 23828
rect 34188 23548 34244 23604
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35644 24556 35700 24612
rect 35756 23938 35812 23940
rect 35756 23886 35758 23938
rect 35758 23886 35810 23938
rect 35810 23886 35812 23938
rect 35756 23884 35812 23886
rect 35252 23772 35308 23828
rect 34972 23436 35028 23492
rect 34412 23378 34468 23380
rect 34412 23326 34414 23378
rect 34414 23326 34466 23378
rect 34466 23326 34468 23378
rect 34412 23324 34468 23326
rect 34300 23154 34356 23156
rect 34300 23102 34302 23154
rect 34302 23102 34354 23154
rect 34354 23102 34356 23154
rect 34300 23100 34356 23102
rect 34524 22988 34580 23044
rect 34300 21756 34356 21812
rect 34188 20972 34244 21028
rect 33628 20802 33684 20804
rect 33628 20750 33630 20802
rect 33630 20750 33682 20802
rect 33682 20750 33684 20802
rect 33628 20748 33684 20750
rect 33740 20076 33796 20132
rect 34076 20636 34132 20692
rect 33964 20188 34020 20244
rect 34300 20076 34356 20132
rect 33180 17948 33236 18004
rect 33068 17612 33124 17668
rect 32396 17052 32452 17108
rect 31836 16268 31892 16324
rect 32060 15932 32116 15988
rect 32396 15484 32452 15540
rect 32172 15260 32228 15316
rect 31836 14924 31892 14980
rect 31724 14364 31780 14420
rect 31836 14700 31892 14756
rect 31948 14588 32004 14644
rect 31724 13634 31780 13636
rect 31724 13582 31726 13634
rect 31726 13582 31778 13634
rect 31778 13582 31780 13634
rect 31724 13580 31780 13582
rect 32284 13580 32340 13636
rect 31948 13074 32004 13076
rect 31948 13022 31950 13074
rect 31950 13022 32002 13074
rect 32002 13022 32004 13074
rect 31948 13020 32004 13022
rect 31724 12236 31780 12292
rect 32620 17388 32676 17444
rect 32956 17442 33012 17444
rect 32956 17390 32958 17442
rect 32958 17390 33010 17442
rect 33010 17390 33012 17442
rect 32956 17388 33012 17390
rect 33180 16940 33236 16996
rect 33292 17500 33348 17556
rect 32956 16380 33012 16436
rect 33180 15314 33236 15316
rect 33180 15262 33182 15314
rect 33182 15262 33234 15314
rect 33234 15262 33236 15314
rect 33180 15260 33236 15262
rect 33852 18226 33908 18228
rect 33852 18174 33854 18226
rect 33854 18174 33906 18226
rect 33906 18174 33908 18226
rect 33852 18172 33908 18174
rect 33740 17778 33796 17780
rect 33740 17726 33742 17778
rect 33742 17726 33794 17778
rect 33794 17726 33796 17778
rect 33740 17724 33796 17726
rect 33404 17388 33460 17444
rect 33628 17442 33684 17444
rect 33628 17390 33630 17442
rect 33630 17390 33682 17442
rect 33682 17390 33684 17442
rect 33628 17388 33684 17390
rect 33404 17106 33460 17108
rect 33404 17054 33406 17106
rect 33406 17054 33458 17106
rect 33458 17054 33460 17106
rect 33404 17052 33460 17054
rect 33404 16098 33460 16100
rect 33404 16046 33406 16098
rect 33406 16046 33458 16098
rect 33458 16046 33460 16098
rect 33404 16044 33460 16046
rect 33740 16380 33796 16436
rect 34412 19964 34468 20020
rect 34300 19234 34356 19236
rect 34300 19182 34302 19234
rect 34302 19182 34354 19234
rect 34354 19182 34356 19234
rect 34300 19180 34356 19182
rect 35420 23436 35476 23492
rect 35644 23548 35700 23604
rect 35196 22988 35252 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 37324 25282 37380 25284
rect 37324 25230 37326 25282
rect 37326 25230 37378 25282
rect 37378 25230 37380 25282
rect 37324 25228 37380 25230
rect 36428 24610 36484 24612
rect 36428 24558 36430 24610
rect 36430 24558 36482 24610
rect 36482 24558 36484 24610
rect 36428 24556 36484 24558
rect 36204 24108 36260 24164
rect 36204 23938 36260 23940
rect 36204 23886 36206 23938
rect 36206 23886 36258 23938
rect 36258 23886 36260 23938
rect 36204 23884 36260 23886
rect 35868 23212 35924 23268
rect 36204 23436 36260 23492
rect 36204 22652 36260 22708
rect 35084 22428 35140 22484
rect 34748 21698 34804 21700
rect 34748 21646 34750 21698
rect 34750 21646 34802 21698
rect 34802 21646 34804 21698
rect 34748 21644 34804 21646
rect 37100 24556 37156 24612
rect 36988 24108 37044 24164
rect 36764 23884 36820 23940
rect 36876 23548 36932 23604
rect 35420 22146 35476 22148
rect 35420 22094 35422 22146
rect 35422 22094 35474 22146
rect 35474 22094 35476 22146
rect 35420 22092 35476 22094
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34636 20076 34692 20132
rect 34524 18674 34580 18676
rect 34524 18622 34526 18674
rect 34526 18622 34578 18674
rect 34578 18622 34580 18674
rect 34524 18620 34580 18622
rect 35084 20690 35140 20692
rect 35084 20638 35086 20690
rect 35086 20638 35138 20690
rect 35138 20638 35140 20690
rect 35084 20636 35140 20638
rect 35980 21756 36036 21812
rect 36876 21698 36932 21700
rect 36876 21646 36878 21698
rect 36878 21646 36930 21698
rect 36930 21646 36932 21698
rect 36876 21644 36932 21646
rect 35868 20802 35924 20804
rect 35868 20750 35870 20802
rect 35870 20750 35922 20802
rect 35922 20750 35924 20802
rect 35868 20748 35924 20750
rect 35420 19906 35476 19908
rect 35420 19854 35422 19906
rect 35422 19854 35474 19906
rect 35474 19854 35476 19906
rect 35420 19852 35476 19854
rect 35644 19740 35700 19796
rect 36092 20690 36148 20692
rect 36092 20638 36094 20690
rect 36094 20638 36146 20690
rect 36146 20638 36148 20690
rect 36092 20636 36148 20638
rect 35868 20130 35924 20132
rect 35868 20078 35870 20130
rect 35870 20078 35922 20130
rect 35922 20078 35924 20130
rect 35868 20076 35924 20078
rect 35756 19964 35812 20020
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 37100 23548 37156 23604
rect 38780 26514 38836 26516
rect 38780 26462 38782 26514
rect 38782 26462 38834 26514
rect 38834 26462 38836 26514
rect 38780 26460 38836 26462
rect 36988 20914 37044 20916
rect 36988 20862 36990 20914
rect 36990 20862 37042 20914
rect 37042 20862 37044 20914
rect 36988 20860 37044 20862
rect 38220 26348 38276 26404
rect 37212 21308 37268 21364
rect 37548 22764 37604 22820
rect 37772 23548 37828 23604
rect 38668 26012 38724 26068
rect 38780 23938 38836 23940
rect 38780 23886 38782 23938
rect 38782 23886 38834 23938
rect 38834 23886 38836 23938
rect 38780 23884 38836 23886
rect 38556 23548 38612 23604
rect 37996 23266 38052 23268
rect 37996 23214 37998 23266
rect 37998 23214 38050 23266
rect 38050 23214 38052 23266
rect 37996 23212 38052 23214
rect 38332 22988 38388 23044
rect 38220 22764 38276 22820
rect 38108 22482 38164 22484
rect 38108 22430 38110 22482
rect 38110 22430 38162 22482
rect 38162 22430 38164 22482
rect 38108 22428 38164 22430
rect 37660 21980 37716 22036
rect 38108 21980 38164 22036
rect 36540 20130 36596 20132
rect 36540 20078 36542 20130
rect 36542 20078 36594 20130
rect 36594 20078 36596 20130
rect 36540 20076 36596 20078
rect 36204 19964 36260 20020
rect 35868 19404 35924 19460
rect 36316 19404 36372 19460
rect 34860 18620 34916 18676
rect 35196 18396 35252 18452
rect 35196 18226 35252 18228
rect 35196 18174 35198 18226
rect 35198 18174 35250 18226
rect 35250 18174 35252 18226
rect 35196 18172 35252 18174
rect 34636 18060 34692 18116
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35756 18620 35812 18676
rect 34524 17724 34580 17780
rect 34748 17554 34804 17556
rect 34748 17502 34750 17554
rect 34750 17502 34802 17554
rect 34802 17502 34804 17554
rect 34748 17500 34804 17502
rect 35084 17666 35140 17668
rect 35084 17614 35086 17666
rect 35086 17614 35138 17666
rect 35138 17614 35140 17666
rect 35084 17612 35140 17614
rect 34188 17164 34244 17220
rect 34300 17052 34356 17108
rect 34412 16994 34468 16996
rect 34412 16942 34414 16994
rect 34414 16942 34466 16994
rect 34466 16942 34468 16994
rect 34412 16940 34468 16942
rect 34412 16716 34468 16772
rect 33740 15426 33796 15428
rect 33740 15374 33742 15426
rect 33742 15374 33794 15426
rect 33794 15374 33796 15426
rect 33740 15372 33796 15374
rect 33628 15260 33684 15316
rect 32508 13692 32564 13748
rect 32172 11564 32228 11620
rect 31724 11228 31780 11284
rect 31836 11170 31892 11172
rect 31836 11118 31838 11170
rect 31838 11118 31890 11170
rect 31890 11118 31892 11170
rect 31836 11116 31892 11118
rect 31612 10892 31668 10948
rect 31612 10722 31668 10724
rect 31612 10670 31614 10722
rect 31614 10670 31666 10722
rect 31666 10670 31668 10722
rect 31612 10668 31668 10670
rect 31500 9884 31556 9940
rect 32284 10444 32340 10500
rect 32956 14364 33012 14420
rect 32732 13580 32788 13636
rect 32620 10444 32676 10500
rect 31052 7756 31108 7812
rect 31836 8876 31892 8932
rect 30604 7196 30660 7252
rect 30604 6018 30660 6020
rect 30604 5966 30606 6018
rect 30606 5966 30658 6018
rect 30658 5966 30660 6018
rect 30604 5964 30660 5966
rect 30156 4172 30212 4228
rect 29708 3836 29764 3892
rect 28476 3500 28532 3556
rect 31500 6412 31556 6468
rect 31164 5906 31220 5908
rect 31164 5854 31166 5906
rect 31166 5854 31218 5906
rect 31218 5854 31220 5906
rect 31164 5852 31220 5854
rect 31276 5404 31332 5460
rect 30940 4732 30996 4788
rect 30828 3836 30884 3892
rect 31500 5292 31556 5348
rect 31836 8428 31892 8484
rect 31612 5180 31668 5236
rect 31724 5740 31780 5796
rect 32732 12684 32788 12740
rect 32508 10220 32564 10276
rect 32396 9100 32452 9156
rect 32508 7980 32564 8036
rect 32284 6690 32340 6692
rect 32284 6638 32286 6690
rect 32286 6638 32338 6690
rect 32338 6638 32340 6690
rect 32284 6636 32340 6638
rect 32172 6524 32228 6580
rect 32172 6018 32228 6020
rect 32172 5966 32174 6018
rect 32174 5966 32226 6018
rect 32226 5966 32228 6018
rect 32172 5964 32228 5966
rect 31948 5906 32004 5908
rect 31948 5854 31950 5906
rect 31950 5854 32002 5906
rect 32002 5854 32004 5906
rect 31948 5852 32004 5854
rect 31836 5628 31892 5684
rect 32060 5292 32116 5348
rect 32396 5122 32452 5124
rect 32396 5070 32398 5122
rect 32398 5070 32450 5122
rect 32450 5070 32452 5122
rect 32396 5068 32452 5070
rect 32172 4956 32228 5012
rect 32172 4226 32228 4228
rect 32172 4174 32174 4226
rect 32174 4174 32226 4226
rect 32226 4174 32228 4226
rect 32172 4172 32228 4174
rect 31612 3554 31668 3556
rect 31612 3502 31614 3554
rect 31614 3502 31666 3554
rect 31666 3502 31668 3554
rect 31612 3500 31668 3502
rect 29484 3442 29540 3444
rect 29484 3390 29486 3442
rect 29486 3390 29538 3442
rect 29538 3390 29540 3442
rect 29484 3388 29540 3390
rect 32396 3442 32452 3444
rect 32396 3390 32398 3442
rect 32398 3390 32450 3442
rect 32450 3390 32452 3442
rect 32396 3388 32452 3390
rect 29484 2828 29540 2884
rect 33180 13634 33236 13636
rect 33180 13582 33182 13634
rect 33182 13582 33234 13634
rect 33234 13582 33236 13634
rect 33180 13580 33236 13582
rect 33404 13356 33460 13412
rect 33516 14924 33572 14980
rect 34076 15372 34132 15428
rect 36876 19852 36932 19908
rect 37212 19740 37268 19796
rect 36540 18956 36596 19012
rect 36652 17836 36708 17892
rect 36540 17778 36596 17780
rect 36540 17726 36542 17778
rect 36542 17726 36594 17778
rect 36594 17726 36596 17778
rect 36540 17724 36596 17726
rect 35980 17276 36036 17332
rect 35308 16716 35364 16772
rect 35196 16604 35252 16660
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35868 15596 35924 15652
rect 34412 15036 34468 15092
rect 34636 15260 34692 15316
rect 34188 14364 34244 14420
rect 33628 13244 33684 13300
rect 34972 15036 35028 15092
rect 34748 14252 34804 14308
rect 33852 13468 33908 13524
rect 34076 13804 34132 13860
rect 33516 12684 33572 12740
rect 33964 12684 34020 12740
rect 33292 10668 33348 10724
rect 33404 10050 33460 10052
rect 33404 9998 33406 10050
rect 33406 9998 33458 10050
rect 33458 9998 33460 10050
rect 33404 9996 33460 9998
rect 32956 9548 33012 9604
rect 33404 9660 33460 9716
rect 33180 9154 33236 9156
rect 33180 9102 33182 9154
rect 33182 9102 33234 9154
rect 33234 9102 33236 9154
rect 33180 9100 33236 9102
rect 33068 9042 33124 9044
rect 33068 8990 33070 9042
rect 33070 8990 33122 9042
rect 33122 8990 33124 9042
rect 33068 8988 33124 8990
rect 32956 8764 33012 8820
rect 34972 14140 35028 14196
rect 34300 13132 34356 13188
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35420 14306 35476 14308
rect 35420 14254 35422 14306
rect 35422 14254 35474 14306
rect 35474 14254 35476 14306
rect 35420 14252 35476 14254
rect 35532 13746 35588 13748
rect 35532 13694 35534 13746
rect 35534 13694 35586 13746
rect 35586 13694 35588 13746
rect 35532 13692 35588 13694
rect 36428 14700 36484 14756
rect 36428 14530 36484 14532
rect 36428 14478 36430 14530
rect 36430 14478 36482 14530
rect 36482 14478 36484 14530
rect 36428 14476 36484 14478
rect 36876 17052 36932 17108
rect 37100 18844 37156 18900
rect 37212 17276 37268 17332
rect 37100 15874 37156 15876
rect 37100 15822 37102 15874
rect 37102 15822 37154 15874
rect 37154 15822 37156 15874
rect 37100 15820 37156 15822
rect 36876 15372 36932 15428
rect 36988 15596 37044 15652
rect 37100 15538 37156 15540
rect 37100 15486 37102 15538
rect 37102 15486 37154 15538
rect 37154 15486 37156 15538
rect 37100 15484 37156 15486
rect 36988 15148 37044 15204
rect 36652 14252 36708 14308
rect 36428 14140 36484 14196
rect 35084 13580 35140 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 12908 35700 12964
rect 34524 11564 34580 11620
rect 34636 12124 34692 12180
rect 35084 12178 35140 12180
rect 35084 12126 35086 12178
rect 35086 12126 35138 12178
rect 35138 12126 35140 12178
rect 35084 12124 35140 12126
rect 33740 8540 33796 8596
rect 33852 8428 33908 8484
rect 34524 10722 34580 10724
rect 34524 10670 34526 10722
rect 34526 10670 34578 10722
rect 34578 10670 34580 10722
rect 34524 10668 34580 10670
rect 34860 11788 34916 11844
rect 34300 9826 34356 9828
rect 34300 9774 34302 9826
rect 34302 9774 34354 9826
rect 34354 9774 34356 9826
rect 34300 9772 34356 9774
rect 34636 8930 34692 8932
rect 34636 8878 34638 8930
rect 34638 8878 34690 8930
rect 34690 8878 34692 8930
rect 34636 8876 34692 8878
rect 34636 8540 34692 8596
rect 32844 7420 32900 7476
rect 32620 5964 32676 6020
rect 33180 6860 33236 6916
rect 33516 6748 33572 6804
rect 33740 7474 33796 7476
rect 33740 7422 33742 7474
rect 33742 7422 33794 7474
rect 33794 7422 33796 7474
rect 33740 7420 33796 7422
rect 33852 6412 33908 6468
rect 33628 5740 33684 5796
rect 34188 7362 34244 7364
rect 34188 7310 34190 7362
rect 34190 7310 34242 7362
rect 34242 7310 34244 7362
rect 34188 7308 34244 7310
rect 34076 6524 34132 6580
rect 33964 5852 34020 5908
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34972 11564 35028 11620
rect 35084 11228 35140 11284
rect 35868 12124 35924 12180
rect 35532 11116 35588 11172
rect 35868 11900 35924 11956
rect 35644 10780 35700 10836
rect 35756 10556 35812 10612
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35084 9772 35140 9828
rect 34972 8034 35028 8036
rect 34972 7982 34974 8034
rect 34974 7982 35026 8034
rect 35026 7982 35028 8034
rect 34972 7980 35028 7982
rect 36092 11452 36148 11508
rect 36316 12738 36372 12740
rect 36316 12686 36318 12738
rect 36318 12686 36370 12738
rect 36370 12686 36372 12738
rect 36316 12684 36372 12686
rect 36428 12178 36484 12180
rect 36428 12126 36430 12178
rect 36430 12126 36482 12178
rect 36482 12126 36484 12178
rect 36428 12124 36484 12126
rect 36204 11170 36260 11172
rect 36204 11118 36206 11170
rect 36206 11118 36258 11170
rect 36258 11118 36260 11170
rect 36204 11116 36260 11118
rect 35868 9884 35924 9940
rect 36204 9602 36260 9604
rect 36204 9550 36206 9602
rect 36206 9550 36258 9602
rect 36258 9550 36260 9602
rect 36204 9548 36260 9550
rect 37100 15036 37156 15092
rect 37100 14418 37156 14420
rect 37100 14366 37102 14418
rect 37102 14366 37154 14418
rect 37154 14366 37156 14418
rect 37100 14364 37156 14366
rect 37100 13634 37156 13636
rect 37100 13582 37102 13634
rect 37102 13582 37154 13634
rect 37154 13582 37156 13634
rect 37100 13580 37156 13582
rect 37100 12850 37156 12852
rect 37100 12798 37102 12850
rect 37102 12798 37154 12850
rect 37154 12798 37156 12850
rect 37100 12796 37156 12798
rect 36876 11452 36932 11508
rect 38444 21362 38500 21364
rect 38444 21310 38446 21362
rect 38446 21310 38498 21362
rect 38498 21310 38500 21362
rect 38444 21308 38500 21310
rect 37996 20802 38052 20804
rect 37996 20750 37998 20802
rect 37998 20750 38050 20802
rect 38050 20750 38052 20802
rect 37996 20748 38052 20750
rect 37436 20130 37492 20132
rect 37436 20078 37438 20130
rect 37438 20078 37490 20130
rect 37490 20078 37492 20130
rect 37436 20076 37492 20078
rect 37996 20018 38052 20020
rect 37996 19966 37998 20018
rect 37998 19966 38050 20018
rect 38050 19966 38052 20018
rect 37996 19964 38052 19966
rect 37436 18956 37492 19012
rect 37884 18844 37940 18900
rect 37996 18450 38052 18452
rect 37996 18398 37998 18450
rect 37998 18398 38050 18450
rect 38050 18398 38052 18450
rect 37996 18396 38052 18398
rect 37772 18060 37828 18116
rect 37548 17778 37604 17780
rect 37548 17726 37550 17778
rect 37550 17726 37602 17778
rect 37602 17726 37604 17778
rect 37548 17724 37604 17726
rect 37548 16882 37604 16884
rect 37548 16830 37550 16882
rect 37550 16830 37602 16882
rect 37602 16830 37604 16882
rect 37548 16828 37604 16830
rect 37436 15820 37492 15876
rect 37436 15596 37492 15652
rect 37324 15372 37380 15428
rect 37772 16828 37828 16884
rect 38220 20860 38276 20916
rect 38444 19628 38500 19684
rect 38220 18956 38276 19012
rect 43372 29148 43428 29204
rect 41020 28476 41076 28532
rect 39676 26572 39732 26628
rect 40236 27132 40292 27188
rect 39004 25506 39060 25508
rect 39004 25454 39006 25506
rect 39006 25454 39058 25506
rect 39058 25454 39060 25506
rect 39004 25452 39060 25454
rect 41580 28476 41636 28532
rect 42028 28364 42084 28420
rect 41356 27858 41412 27860
rect 41356 27806 41358 27858
rect 41358 27806 41410 27858
rect 41410 27806 41412 27858
rect 41356 27804 41412 27806
rect 41020 27186 41076 27188
rect 41020 27134 41022 27186
rect 41022 27134 41074 27186
rect 41074 27134 41076 27186
rect 41020 27132 41076 27134
rect 42252 27580 42308 27636
rect 41468 27074 41524 27076
rect 41468 27022 41470 27074
rect 41470 27022 41522 27074
rect 41522 27022 41524 27074
rect 41468 27020 41524 27022
rect 39676 26402 39732 26404
rect 39676 26350 39678 26402
rect 39678 26350 39730 26402
rect 39730 26350 39732 26402
rect 39676 26348 39732 26350
rect 39228 26012 39284 26068
rect 41244 25228 41300 25284
rect 40348 23826 40404 23828
rect 40348 23774 40350 23826
rect 40350 23774 40402 23826
rect 40402 23774 40404 23826
rect 40348 23772 40404 23774
rect 40012 23212 40068 23268
rect 39004 23042 39060 23044
rect 39004 22990 39006 23042
rect 39006 22990 39058 23042
rect 39058 22990 39060 23042
rect 39004 22988 39060 22990
rect 39116 22876 39172 22932
rect 39004 22652 39060 22708
rect 39228 22764 39284 22820
rect 39452 21868 39508 21924
rect 39676 22930 39732 22932
rect 39676 22878 39678 22930
rect 39678 22878 39730 22930
rect 39730 22878 39732 22930
rect 39676 22876 39732 22878
rect 39788 22652 39844 22708
rect 40124 23154 40180 23156
rect 40124 23102 40126 23154
rect 40126 23102 40178 23154
rect 40178 23102 40180 23154
rect 40124 23100 40180 23102
rect 40124 22764 40180 22820
rect 38444 18172 38500 18228
rect 38108 17052 38164 17108
rect 37996 16940 38052 16996
rect 37884 15820 37940 15876
rect 37660 15036 37716 15092
rect 37548 14924 37604 14980
rect 38220 15820 38276 15876
rect 38108 15596 38164 15652
rect 38780 17666 38836 17668
rect 38780 17614 38782 17666
rect 38782 17614 38834 17666
rect 38834 17614 38836 17666
rect 38780 17612 38836 17614
rect 38892 17276 38948 17332
rect 38332 15484 38388 15540
rect 38668 17164 38724 17220
rect 38108 14924 38164 14980
rect 37660 14418 37716 14420
rect 37660 14366 37662 14418
rect 37662 14366 37714 14418
rect 37714 14366 37716 14418
rect 37660 14364 37716 14366
rect 37548 13522 37604 13524
rect 37548 13470 37550 13522
rect 37550 13470 37602 13522
rect 37602 13470 37604 13522
rect 37548 13468 37604 13470
rect 37884 14306 37940 14308
rect 37884 14254 37886 14306
rect 37886 14254 37938 14306
rect 37938 14254 37940 14306
rect 37884 14252 37940 14254
rect 37772 13468 37828 13524
rect 37548 13132 37604 13188
rect 37660 12908 37716 12964
rect 37324 12290 37380 12292
rect 37324 12238 37326 12290
rect 37326 12238 37378 12290
rect 37378 12238 37380 12290
rect 37324 12236 37380 12238
rect 37772 11676 37828 11732
rect 37100 10668 37156 10724
rect 37660 10668 37716 10724
rect 36204 8876 36260 8932
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35644 8316 35700 8372
rect 36204 8316 36260 8372
rect 34748 7474 34804 7476
rect 34748 7422 34750 7474
rect 34750 7422 34802 7474
rect 34802 7422 34804 7474
rect 34748 7420 34804 7422
rect 34524 6466 34580 6468
rect 34524 6414 34526 6466
rect 34526 6414 34578 6466
rect 34578 6414 34580 6466
rect 34524 6412 34580 6414
rect 34076 6076 34132 6132
rect 34972 7308 35028 7364
rect 33292 5234 33348 5236
rect 33292 5182 33294 5234
rect 33294 5182 33346 5234
rect 33346 5182 33348 5234
rect 33292 5180 33348 5182
rect 33180 4956 33236 5012
rect 33180 4732 33236 4788
rect 33740 5122 33796 5124
rect 33740 5070 33742 5122
rect 33742 5070 33794 5122
rect 33794 5070 33796 5122
rect 33740 5068 33796 5070
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 6860 35252 6916
rect 35644 7362 35700 7364
rect 35644 7310 35646 7362
rect 35646 7310 35698 7362
rect 35698 7310 35700 7362
rect 35644 7308 35700 7310
rect 35644 6188 35700 6244
rect 35196 6018 35252 6020
rect 35196 5966 35198 6018
rect 35198 5966 35250 6018
rect 35250 5966 35252 6018
rect 35196 5964 35252 5966
rect 36316 8146 36372 8148
rect 36316 8094 36318 8146
rect 36318 8094 36370 8146
rect 36370 8094 36372 8146
rect 36316 8092 36372 8094
rect 37996 11394 38052 11396
rect 37996 11342 37998 11394
rect 37998 11342 38050 11394
rect 38050 11342 38052 11394
rect 37996 11340 38052 11342
rect 37884 11116 37940 11172
rect 37100 9938 37156 9940
rect 37100 9886 37102 9938
rect 37102 9886 37154 9938
rect 37154 9886 37156 9938
rect 37100 9884 37156 9886
rect 36652 7698 36708 7700
rect 36652 7646 36654 7698
rect 36654 7646 36706 7698
rect 36706 7646 36708 7698
rect 36652 7644 36708 7646
rect 36540 7532 36596 7588
rect 36988 8316 37044 8372
rect 37100 9100 37156 9156
rect 37996 9826 38052 9828
rect 37996 9774 37998 9826
rect 37998 9774 38050 9826
rect 38050 9774 38052 9826
rect 37996 9772 38052 9774
rect 38220 12908 38276 12964
rect 38556 15148 38612 15204
rect 38332 14028 38388 14084
rect 38444 14364 38500 14420
rect 38444 13020 38500 13076
rect 39116 17388 39172 17444
rect 39116 16940 39172 16996
rect 38892 16716 38948 16772
rect 38892 15596 38948 15652
rect 39564 18284 39620 18340
rect 40012 19628 40068 19684
rect 39788 18450 39844 18452
rect 39788 18398 39790 18450
rect 39790 18398 39842 18450
rect 39842 18398 39844 18450
rect 39788 18396 39844 18398
rect 39676 18060 39732 18116
rect 39900 17612 39956 17668
rect 39676 17442 39732 17444
rect 39676 17390 39678 17442
rect 39678 17390 39730 17442
rect 39730 17390 39732 17442
rect 39676 17388 39732 17390
rect 39788 17052 39844 17108
rect 39564 16156 39620 16212
rect 38668 14700 38724 14756
rect 38668 13692 38724 13748
rect 38892 13468 38948 13524
rect 38220 12738 38276 12740
rect 38220 12686 38222 12738
rect 38222 12686 38274 12738
rect 38274 12686 38276 12738
rect 38220 12684 38276 12686
rect 38556 12738 38612 12740
rect 38556 12686 38558 12738
rect 38558 12686 38610 12738
rect 38610 12686 38612 12738
rect 38556 12684 38612 12686
rect 38220 12348 38276 12404
rect 39340 14924 39396 14980
rect 39788 14812 39844 14868
rect 39900 14700 39956 14756
rect 40124 16716 40180 16772
rect 42812 28418 42868 28420
rect 42812 28366 42814 28418
rect 42814 28366 42866 28418
rect 42866 28366 42868 28418
rect 42812 28364 42868 28366
rect 43260 27580 43316 27636
rect 45276 29202 45332 29204
rect 45276 29150 45278 29202
rect 45278 29150 45330 29202
rect 45330 29150 45332 29202
rect 45276 29148 45332 29150
rect 44492 28476 44548 28532
rect 45164 28364 45220 28420
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 45052 27634 45108 27636
rect 45052 27582 45054 27634
rect 45054 27582 45106 27634
rect 45106 27582 45108 27634
rect 45052 27580 45108 27582
rect 43596 27132 43652 27188
rect 43596 26908 43652 26964
rect 42364 25564 42420 25620
rect 43148 26236 43204 26292
rect 42364 25340 42420 25396
rect 42028 23714 42084 23716
rect 42028 23662 42030 23714
rect 42030 23662 42082 23714
rect 42082 23662 42084 23714
rect 42028 23660 42084 23662
rect 41020 23266 41076 23268
rect 41020 23214 41022 23266
rect 41022 23214 41074 23266
rect 41074 23214 41076 23266
rect 41020 23212 41076 23214
rect 41804 23266 41860 23268
rect 41804 23214 41806 23266
rect 41806 23214 41858 23266
rect 41858 23214 41860 23266
rect 41804 23212 41860 23214
rect 40908 23154 40964 23156
rect 40908 23102 40910 23154
rect 40910 23102 40962 23154
rect 40962 23102 40964 23154
rect 40908 23100 40964 23102
rect 42140 23042 42196 23044
rect 42140 22990 42142 23042
rect 42142 22990 42194 23042
rect 42194 22990 42196 23042
rect 42140 22988 42196 22990
rect 40796 22652 40852 22708
rect 41020 22764 41076 22820
rect 41916 22764 41972 22820
rect 41132 22092 41188 22148
rect 40460 21420 40516 21476
rect 40572 20690 40628 20692
rect 40572 20638 40574 20690
rect 40574 20638 40626 20690
rect 40626 20638 40628 20690
rect 40572 20636 40628 20638
rect 41244 21474 41300 21476
rect 41244 21422 41246 21474
rect 41246 21422 41298 21474
rect 41298 21422 41300 21474
rect 41244 21420 41300 21422
rect 41468 21420 41524 21476
rect 42588 24780 42644 24836
rect 42364 22764 42420 22820
rect 42140 21756 42196 21812
rect 41916 21308 41972 21364
rect 41580 20636 41636 20692
rect 42140 20636 42196 20692
rect 42252 21420 42308 21476
rect 41692 20412 41748 20468
rect 41804 19906 41860 19908
rect 41804 19854 41806 19906
rect 41806 19854 41858 19906
rect 41858 19854 41860 19906
rect 41804 19852 41860 19854
rect 41020 17724 41076 17780
rect 40348 16716 40404 16772
rect 41132 17554 41188 17556
rect 41132 17502 41134 17554
rect 41134 17502 41186 17554
rect 41186 17502 41188 17554
rect 41132 17500 41188 17502
rect 41244 17388 41300 17444
rect 41468 16828 41524 16884
rect 41356 16716 41412 16772
rect 40908 16604 40964 16660
rect 41804 18396 41860 18452
rect 42140 18956 42196 19012
rect 41916 18284 41972 18340
rect 41804 17500 41860 17556
rect 41692 17388 41748 17444
rect 42028 17442 42084 17444
rect 42028 17390 42030 17442
rect 42030 17390 42082 17442
rect 42082 17390 42084 17442
rect 42028 17388 42084 17390
rect 41916 17276 41972 17332
rect 41804 16770 41860 16772
rect 41804 16718 41806 16770
rect 41806 16718 41858 16770
rect 41858 16718 41860 16770
rect 41804 16716 41860 16718
rect 40348 16268 40404 16324
rect 41244 15202 41300 15204
rect 41244 15150 41246 15202
rect 41246 15150 41298 15202
rect 41298 15150 41300 15202
rect 41244 15148 41300 15150
rect 40236 14924 40292 14980
rect 40124 14364 40180 14420
rect 38780 11676 38836 11732
rect 38444 11506 38500 11508
rect 38444 11454 38446 11506
rect 38446 11454 38498 11506
rect 38498 11454 38500 11506
rect 38444 11452 38500 11454
rect 38108 9100 38164 9156
rect 38332 10668 38388 10724
rect 38556 11170 38612 11172
rect 38556 11118 38558 11170
rect 38558 11118 38610 11170
rect 38610 11118 38612 11170
rect 38556 11116 38612 11118
rect 38556 9938 38612 9940
rect 38556 9886 38558 9938
rect 38558 9886 38610 9938
rect 38610 9886 38612 9938
rect 38556 9884 38612 9886
rect 38892 9884 38948 9940
rect 39452 12684 39508 12740
rect 39564 12178 39620 12180
rect 39564 12126 39566 12178
rect 39566 12126 39618 12178
rect 39618 12126 39620 12178
rect 39564 12124 39620 12126
rect 38780 9154 38836 9156
rect 38780 9102 38782 9154
rect 38782 9102 38834 9154
rect 38834 9102 38836 9154
rect 38780 9100 38836 9102
rect 37884 8316 37940 8372
rect 37212 8146 37268 8148
rect 37212 8094 37214 8146
rect 37214 8094 37266 8146
rect 37266 8094 37268 8146
rect 37212 8092 37268 8094
rect 38444 8146 38500 8148
rect 38444 8094 38446 8146
rect 38446 8094 38498 8146
rect 38498 8094 38500 8146
rect 38444 8092 38500 8094
rect 37548 7644 37604 7700
rect 36316 6188 36372 6244
rect 36540 6524 36596 6580
rect 36092 5628 36148 5684
rect 37100 7308 37156 7364
rect 38668 7474 38724 7476
rect 38668 7422 38670 7474
rect 38670 7422 38722 7474
rect 38722 7422 38724 7474
rect 38668 7420 38724 7422
rect 37996 7362 38052 7364
rect 37996 7310 37998 7362
rect 37998 7310 38050 7362
rect 38050 7310 38052 7362
rect 37996 7308 38052 7310
rect 37548 7196 37604 7252
rect 38332 7250 38388 7252
rect 38332 7198 38334 7250
rect 38334 7198 38386 7250
rect 38386 7198 38388 7250
rect 38332 7196 38388 7198
rect 37996 6690 38052 6692
rect 37996 6638 37998 6690
rect 37998 6638 38050 6690
rect 38050 6638 38052 6690
rect 37996 6636 38052 6638
rect 38444 6578 38500 6580
rect 38444 6526 38446 6578
rect 38446 6526 38498 6578
rect 38498 6526 38500 6578
rect 38444 6524 38500 6526
rect 37324 6188 37380 6244
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35420 5292 35476 5348
rect 34524 4562 34580 4564
rect 34524 4510 34526 4562
rect 34526 4510 34578 4562
rect 34578 4510 34580 4562
rect 34524 4508 34580 4510
rect 35196 3946 35252 3948
rect 33180 3836 33236 3892
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34076 3666 34132 3668
rect 34076 3614 34078 3666
rect 34078 3614 34130 3666
rect 34130 3614 34132 3666
rect 34076 3612 34132 3614
rect 32732 3330 32788 3332
rect 32732 3278 32734 3330
rect 32734 3278 32786 3330
rect 32786 3278 32788 3330
rect 32732 3276 32788 3278
rect 38892 5628 38948 5684
rect 38780 3052 38836 3108
rect 36876 2604 36932 2660
rect 32508 2380 32564 2436
rect 26908 1596 26964 1652
rect 40012 14028 40068 14084
rect 39900 13746 39956 13748
rect 39900 13694 39902 13746
rect 39902 13694 39954 13746
rect 39954 13694 39956 13746
rect 39900 13692 39956 13694
rect 41020 14812 41076 14868
rect 40460 12908 40516 12964
rect 40012 12796 40068 12852
rect 39900 12348 39956 12404
rect 40124 12684 40180 12740
rect 39900 10780 39956 10836
rect 39340 9714 39396 9716
rect 39340 9662 39342 9714
rect 39342 9662 39394 9714
rect 39394 9662 39396 9714
rect 39340 9660 39396 9662
rect 39564 9996 39620 10052
rect 40684 13020 40740 13076
rect 40908 13580 40964 13636
rect 41020 13468 41076 13524
rect 40796 12572 40852 12628
rect 41244 12460 41300 12516
rect 40684 12124 40740 12180
rect 39116 7420 39172 7476
rect 39340 8988 39396 9044
rect 39900 8204 39956 8260
rect 40236 6748 40292 6804
rect 40572 9714 40628 9716
rect 40572 9662 40574 9714
rect 40574 9662 40626 9714
rect 40626 9662 40628 9714
rect 40572 9660 40628 9662
rect 41468 15260 41524 15316
rect 41916 16604 41972 16660
rect 42140 16828 42196 16884
rect 42028 16492 42084 16548
rect 42476 21308 42532 21364
rect 42700 23660 42756 23716
rect 43708 26290 43764 26292
rect 43708 26238 43710 26290
rect 43710 26238 43762 26290
rect 43762 26238 43764 26290
rect 43708 26236 43764 26238
rect 42812 23212 42868 23268
rect 42812 21868 42868 21924
rect 42812 21586 42868 21588
rect 42812 21534 42814 21586
rect 42814 21534 42866 21586
rect 42866 21534 42868 21586
rect 42812 21532 42868 21534
rect 42812 20412 42868 20468
rect 45164 25452 45220 25508
rect 43372 25394 43428 25396
rect 43372 25342 43374 25394
rect 43374 25342 43426 25394
rect 43426 25342 43428 25394
rect 43372 25340 43428 25342
rect 43372 24834 43428 24836
rect 43372 24782 43374 24834
rect 43374 24782 43426 24834
rect 43426 24782 43428 24834
rect 43372 24780 43428 24782
rect 43148 24162 43204 24164
rect 43148 24110 43150 24162
rect 43150 24110 43202 24162
rect 43202 24110 43204 24162
rect 43148 24108 43204 24110
rect 43484 24668 43540 24724
rect 44716 24722 44772 24724
rect 44716 24670 44718 24722
rect 44718 24670 44770 24722
rect 44770 24670 44772 24722
rect 44716 24668 44772 24670
rect 44380 24610 44436 24612
rect 44380 24558 44382 24610
rect 44382 24558 44434 24610
rect 44434 24558 44436 24610
rect 44380 24556 44436 24558
rect 43148 23212 43204 23268
rect 43036 21868 43092 21924
rect 42588 18396 42644 18452
rect 42924 18284 42980 18340
rect 42588 18172 42644 18228
rect 42812 17890 42868 17892
rect 42812 17838 42814 17890
rect 42814 17838 42866 17890
rect 42866 17838 42868 17890
rect 42812 17836 42868 17838
rect 42700 17554 42756 17556
rect 42700 17502 42702 17554
rect 42702 17502 42754 17554
rect 42754 17502 42756 17554
rect 42700 17500 42756 17502
rect 42364 16492 42420 16548
rect 42476 16156 42532 16212
rect 42028 15426 42084 15428
rect 42028 15374 42030 15426
rect 42030 15374 42082 15426
rect 42082 15374 42084 15426
rect 42028 15372 42084 15374
rect 42028 15036 42084 15092
rect 42028 13468 42084 13524
rect 41468 12850 41524 12852
rect 41468 12798 41470 12850
rect 41470 12798 41522 12850
rect 41522 12798 41524 12850
rect 41468 12796 41524 12798
rect 41356 10780 41412 10836
rect 41468 10556 41524 10612
rect 41020 9996 41076 10052
rect 40684 9100 40740 9156
rect 41244 8764 41300 8820
rect 40572 8258 40628 8260
rect 40572 8206 40574 8258
rect 40574 8206 40626 8258
rect 40626 8206 40628 8258
rect 40572 8204 40628 8206
rect 41692 12738 41748 12740
rect 41692 12686 41694 12738
rect 41694 12686 41746 12738
rect 41746 12686 41748 12738
rect 41692 12684 41748 12686
rect 42476 15372 42532 15428
rect 42364 13074 42420 13076
rect 42364 13022 42366 13074
rect 42366 13022 42418 13074
rect 42418 13022 42420 13074
rect 42364 13020 42420 13022
rect 42476 12460 42532 12516
rect 42364 12012 42420 12068
rect 42252 11900 42308 11956
rect 41692 10834 41748 10836
rect 41692 10782 41694 10834
rect 41694 10782 41746 10834
rect 41746 10782 41748 10834
rect 41692 10780 41748 10782
rect 42028 10556 42084 10612
rect 42252 10444 42308 10500
rect 41804 9996 41860 10052
rect 42812 17164 42868 17220
rect 43036 16044 43092 16100
rect 42700 15874 42756 15876
rect 42700 15822 42702 15874
rect 42702 15822 42754 15874
rect 42754 15822 42756 15874
rect 42700 15820 42756 15822
rect 42924 15260 42980 15316
rect 42812 14306 42868 14308
rect 42812 14254 42814 14306
rect 42814 14254 42866 14306
rect 42866 14254 42868 14306
rect 42812 14252 42868 14254
rect 44268 23436 44324 23492
rect 43372 22146 43428 22148
rect 43372 22094 43374 22146
rect 43374 22094 43426 22146
rect 43426 22094 43428 22146
rect 43372 22092 43428 22094
rect 43596 23100 43652 23156
rect 43596 21868 43652 21924
rect 43708 22428 43764 22484
rect 44156 23154 44212 23156
rect 44156 23102 44158 23154
rect 44158 23102 44210 23154
rect 44210 23102 44212 23154
rect 44156 23100 44212 23102
rect 44492 22540 44548 22596
rect 43484 21586 43540 21588
rect 43484 21534 43486 21586
rect 43486 21534 43538 21586
rect 43538 21534 43540 21586
rect 43484 21532 43540 21534
rect 43820 22370 43876 22372
rect 43820 22318 43822 22370
rect 43822 22318 43874 22370
rect 43874 22318 43876 22370
rect 43820 22316 43876 22318
rect 43932 22146 43988 22148
rect 43932 22094 43934 22146
rect 43934 22094 43986 22146
rect 43986 22094 43988 22146
rect 43932 22092 43988 22094
rect 44156 21868 44212 21924
rect 46396 27356 46452 27412
rect 49644 27858 49700 27860
rect 49644 27806 49646 27858
rect 49646 27806 49698 27858
rect 49698 27806 49700 27858
rect 49644 27804 49700 27806
rect 47964 27746 48020 27748
rect 47964 27694 47966 27746
rect 47966 27694 48018 27746
rect 48018 27694 48020 27746
rect 47964 27692 48020 27694
rect 45612 26908 45668 26964
rect 45836 26962 45892 26964
rect 45836 26910 45838 26962
rect 45838 26910 45890 26962
rect 45890 26910 45892 26962
rect 45836 26908 45892 26910
rect 46508 26908 46564 26964
rect 46844 27356 46900 27412
rect 47404 27356 47460 27412
rect 49420 27356 49476 27412
rect 49532 27692 49588 27748
rect 49084 27298 49140 27300
rect 49084 27246 49086 27298
rect 49086 27246 49138 27298
rect 49138 27246 49140 27298
rect 49084 27244 49140 27246
rect 48748 26962 48804 26964
rect 48748 26910 48750 26962
rect 48750 26910 48802 26962
rect 48802 26910 48804 26962
rect 48748 26908 48804 26910
rect 44940 23436 44996 23492
rect 45388 23324 45444 23380
rect 45388 22540 45444 22596
rect 45500 22092 45556 22148
rect 44940 21868 44996 21924
rect 44828 21756 44884 21812
rect 43932 19292 43988 19348
rect 43596 18620 43652 18676
rect 43372 18396 43428 18452
rect 44156 18284 44212 18340
rect 44604 18284 44660 18340
rect 43260 17836 43316 17892
rect 43596 16044 43652 16100
rect 43372 15932 43428 15988
rect 43148 14418 43204 14420
rect 43148 14366 43150 14418
rect 43150 14366 43202 14418
rect 43202 14366 43204 14418
rect 43148 14364 43204 14366
rect 42924 13580 42980 13636
rect 42812 13468 42868 13524
rect 42812 12012 42868 12068
rect 43148 11900 43204 11956
rect 43932 16098 43988 16100
rect 43932 16046 43934 16098
rect 43934 16046 43986 16098
rect 43986 16046 43988 16098
rect 43932 16044 43988 16046
rect 44156 16044 44212 16100
rect 45388 20524 45444 20580
rect 45276 19964 45332 20020
rect 44828 18508 44884 18564
rect 45164 17554 45220 17556
rect 45164 17502 45166 17554
rect 45166 17502 45218 17554
rect 45218 17502 45220 17554
rect 45164 17500 45220 17502
rect 45052 16716 45108 16772
rect 45500 19964 45556 20020
rect 45724 18620 45780 18676
rect 46508 26124 46564 26180
rect 46284 25506 46340 25508
rect 46284 25454 46286 25506
rect 46286 25454 46338 25506
rect 46338 25454 46340 25506
rect 46284 25452 46340 25454
rect 49868 27746 49924 27748
rect 49868 27694 49870 27746
rect 49870 27694 49922 27746
rect 49922 27694 49924 27746
rect 49868 27692 49924 27694
rect 50428 27692 50484 27748
rect 50316 27634 50372 27636
rect 50316 27582 50318 27634
rect 50318 27582 50370 27634
rect 50370 27582 50372 27634
rect 50316 27580 50372 27582
rect 49980 27356 50036 27412
rect 49644 27244 49700 27300
rect 51100 27858 51156 27860
rect 51100 27806 51102 27858
rect 51102 27806 51154 27858
rect 51154 27806 51156 27858
rect 51100 27804 51156 27806
rect 51996 27858 52052 27860
rect 51996 27806 51998 27858
rect 51998 27806 52050 27858
rect 52050 27806 52052 27858
rect 51996 27804 52052 27806
rect 50876 27356 50932 27412
rect 51660 27634 51716 27636
rect 51660 27582 51662 27634
rect 51662 27582 51714 27634
rect 51714 27582 51716 27634
rect 51660 27580 51716 27582
rect 51772 27074 51828 27076
rect 51772 27022 51774 27074
rect 51774 27022 51826 27074
rect 51826 27022 51828 27074
rect 51772 27020 51828 27022
rect 49756 26402 49812 26404
rect 49756 26350 49758 26402
rect 49758 26350 49810 26402
rect 49810 26350 49812 26402
rect 49756 26348 49812 26350
rect 46956 26178 47012 26180
rect 46956 26126 46958 26178
rect 46958 26126 47010 26178
rect 47010 26126 47012 26178
rect 46956 26124 47012 26126
rect 47180 25618 47236 25620
rect 47180 25566 47182 25618
rect 47182 25566 47234 25618
rect 47234 25566 47236 25618
rect 47180 25564 47236 25566
rect 50876 26908 50932 26964
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50316 26402 50372 26404
rect 50316 26350 50318 26402
rect 50318 26350 50370 26402
rect 50370 26350 50372 26402
rect 50316 26348 50372 26350
rect 50092 26236 50148 26292
rect 49084 25564 49140 25620
rect 46844 25452 46900 25508
rect 48860 25452 48916 25508
rect 46508 25228 46564 25284
rect 46956 25228 47012 25284
rect 46284 24722 46340 24724
rect 46284 24670 46286 24722
rect 46286 24670 46338 24722
rect 46338 24670 46340 24722
rect 46284 24668 46340 24670
rect 46060 21980 46116 22036
rect 45948 21868 46004 21924
rect 45500 17666 45556 17668
rect 45500 17614 45502 17666
rect 45502 17614 45554 17666
rect 45554 17614 45556 17666
rect 45500 17612 45556 17614
rect 45500 16716 45556 16772
rect 44828 15986 44884 15988
rect 44828 15934 44830 15986
rect 44830 15934 44882 15986
rect 44882 15934 44884 15986
rect 44828 15932 44884 15934
rect 45164 15708 45220 15764
rect 46172 21308 46228 21364
rect 46844 24162 46900 24164
rect 46844 24110 46846 24162
rect 46846 24110 46898 24162
rect 46898 24110 46900 24162
rect 46844 24108 46900 24110
rect 50988 26290 51044 26292
rect 50988 26238 50990 26290
rect 50990 26238 51042 26290
rect 51042 26238 51044 26290
rect 50988 26236 51044 26238
rect 51436 26236 51492 26292
rect 50540 25900 50596 25956
rect 50204 25452 50260 25508
rect 50652 25506 50708 25508
rect 50652 25454 50654 25506
rect 50654 25454 50706 25506
rect 50706 25454 50708 25506
rect 50652 25452 50708 25454
rect 50876 25900 50932 25956
rect 52892 27858 52948 27860
rect 52892 27806 52894 27858
rect 52894 27806 52946 27858
rect 52946 27806 52948 27858
rect 52892 27804 52948 27806
rect 51996 27020 52052 27076
rect 57932 27580 57988 27636
rect 54236 27020 54292 27076
rect 55580 27074 55636 27076
rect 55580 27022 55582 27074
rect 55582 27022 55634 27074
rect 55634 27022 55636 27074
rect 55580 27020 55636 27022
rect 52556 26908 52612 26964
rect 52332 26290 52388 26292
rect 52332 26238 52334 26290
rect 52334 26238 52386 26290
rect 52386 26238 52388 26290
rect 52332 26236 52388 26238
rect 52892 26236 52948 26292
rect 53676 26290 53732 26292
rect 53676 26238 53678 26290
rect 53678 26238 53730 26290
rect 53730 26238 53732 26290
rect 53676 26236 53732 26238
rect 51660 25564 51716 25620
rect 52668 25618 52724 25620
rect 52668 25566 52670 25618
rect 52670 25566 52722 25618
rect 52722 25566 52724 25618
rect 52668 25564 52724 25566
rect 50764 25228 50820 25284
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 47068 24722 47124 24724
rect 47068 24670 47070 24722
rect 47070 24670 47122 24722
rect 47122 24670 47124 24722
rect 47068 24668 47124 24670
rect 47964 24668 48020 24724
rect 47180 23884 47236 23940
rect 46172 20524 46228 20580
rect 46396 20636 46452 20692
rect 46844 21586 46900 21588
rect 46844 21534 46846 21586
rect 46846 21534 46898 21586
rect 46898 21534 46900 21586
rect 46844 21532 46900 21534
rect 46620 20188 46676 20244
rect 46844 20076 46900 20132
rect 46620 19234 46676 19236
rect 46620 19182 46622 19234
rect 46622 19182 46674 19234
rect 46674 19182 46676 19234
rect 46620 19180 46676 19182
rect 46060 19010 46116 19012
rect 46060 18958 46062 19010
rect 46062 18958 46114 19010
rect 46114 18958 46116 19010
rect 46060 18956 46116 18958
rect 46284 19010 46340 19012
rect 46284 18958 46286 19010
rect 46286 18958 46338 19010
rect 46338 18958 46340 19010
rect 46284 18956 46340 18958
rect 46060 16770 46116 16772
rect 46060 16718 46062 16770
rect 46062 16718 46114 16770
rect 46114 16718 46116 16770
rect 46060 16716 46116 16718
rect 43484 14306 43540 14308
rect 43484 14254 43486 14306
rect 43486 14254 43538 14306
rect 43538 14254 43540 14306
rect 43484 14252 43540 14254
rect 43372 12908 43428 12964
rect 43260 11452 43316 11508
rect 42812 11004 42868 11060
rect 42812 10444 42868 10500
rect 40908 6690 40964 6692
rect 40908 6638 40910 6690
rect 40910 6638 40962 6690
rect 40962 6638 40964 6690
rect 40908 6636 40964 6638
rect 41356 6690 41412 6692
rect 41356 6638 41358 6690
rect 41358 6638 41410 6690
rect 41410 6638 41412 6690
rect 41356 6636 41412 6638
rect 40348 6412 40404 6468
rect 42028 9154 42084 9156
rect 42028 9102 42030 9154
rect 42030 9102 42082 9154
rect 42082 9102 42084 9154
rect 42028 9100 42084 9102
rect 41916 7250 41972 7252
rect 41916 7198 41918 7250
rect 41918 7198 41970 7250
rect 41970 7198 41972 7250
rect 41916 7196 41972 7198
rect 41916 6578 41972 6580
rect 41916 6526 41918 6578
rect 41918 6526 41970 6578
rect 41970 6526 41972 6578
rect 41916 6524 41972 6526
rect 39452 5682 39508 5684
rect 39452 5630 39454 5682
rect 39454 5630 39506 5682
rect 39506 5630 39508 5682
rect 39452 5628 39508 5630
rect 39788 5122 39844 5124
rect 39788 5070 39790 5122
rect 39790 5070 39842 5122
rect 39842 5070 39844 5122
rect 39788 5068 39844 5070
rect 41132 5234 41188 5236
rect 41132 5182 41134 5234
rect 41134 5182 41186 5234
rect 41186 5182 41188 5234
rect 41132 5180 41188 5182
rect 39676 4956 39732 5012
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 43372 10892 43428 10948
rect 43260 10610 43316 10612
rect 43260 10558 43262 10610
rect 43262 10558 43314 10610
rect 43314 10558 43316 10610
rect 43260 10556 43316 10558
rect 43932 12908 43988 12964
rect 43820 12124 43876 12180
rect 43484 9996 43540 10052
rect 42924 9602 42980 9604
rect 42924 9550 42926 9602
rect 42926 9550 42978 9602
rect 42978 9550 42980 9602
rect 42924 9548 42980 9550
rect 42812 9100 42868 9156
rect 43484 9602 43540 9604
rect 43484 9550 43486 9602
rect 43486 9550 43538 9602
rect 43538 9550 43540 9602
rect 43484 9548 43540 9550
rect 45388 13746 45444 13748
rect 45388 13694 45390 13746
rect 45390 13694 45442 13746
rect 45442 13694 45444 13746
rect 45388 13692 45444 13694
rect 45500 14476 45556 14532
rect 44268 12962 44324 12964
rect 44268 12910 44270 12962
rect 44270 12910 44322 12962
rect 44322 12910 44324 12962
rect 44268 12908 44324 12910
rect 45388 12178 45444 12180
rect 45388 12126 45390 12178
rect 45390 12126 45442 12178
rect 45442 12126 45444 12178
rect 45388 12124 45444 12126
rect 46172 16098 46228 16100
rect 46172 16046 46174 16098
rect 46174 16046 46226 16098
rect 46226 16046 46228 16098
rect 46172 16044 46228 16046
rect 45948 14812 46004 14868
rect 46508 15708 46564 15764
rect 46956 19852 47012 19908
rect 48188 23884 48244 23940
rect 48972 24722 49028 24724
rect 48972 24670 48974 24722
rect 48974 24670 49026 24722
rect 49026 24670 49028 24722
rect 48972 24668 49028 24670
rect 48748 23884 48804 23940
rect 49308 24556 49364 24612
rect 47964 23548 48020 23604
rect 47628 23212 47684 23268
rect 47292 22988 47348 23044
rect 47292 22482 47348 22484
rect 47292 22430 47294 22482
rect 47294 22430 47346 22482
rect 47346 22430 47348 22482
rect 47292 22428 47348 22430
rect 47404 21980 47460 22036
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 51436 23436 51492 23492
rect 50204 23324 50260 23380
rect 51100 23324 51156 23380
rect 52780 23436 52836 23492
rect 51884 23324 51940 23380
rect 51212 23266 51268 23268
rect 51212 23214 51214 23266
rect 51214 23214 51266 23266
rect 51266 23214 51268 23266
rect 51212 23212 51268 23214
rect 51660 23266 51716 23268
rect 51660 23214 51662 23266
rect 51662 23214 51714 23266
rect 51714 23214 51716 23266
rect 51660 23212 51716 23214
rect 52220 23378 52276 23380
rect 52220 23326 52222 23378
rect 52222 23326 52274 23378
rect 52274 23326 52276 23378
rect 52220 23324 52276 23326
rect 52892 23324 52948 23380
rect 47964 22594 48020 22596
rect 47964 22542 47966 22594
rect 47966 22542 48018 22594
rect 48018 22542 48020 22594
rect 47964 22540 48020 22542
rect 47740 22428 47796 22484
rect 50876 22428 50932 22484
rect 50204 22370 50260 22372
rect 50204 22318 50206 22370
rect 50206 22318 50258 22370
rect 50258 22318 50260 22370
rect 50204 22316 50260 22318
rect 50652 22092 50708 22148
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 49420 21698 49476 21700
rect 49420 21646 49422 21698
rect 49422 21646 49474 21698
rect 49474 21646 49476 21698
rect 49420 21644 49476 21646
rect 47404 21532 47460 21588
rect 49196 21084 49252 21140
rect 47740 20690 47796 20692
rect 47740 20638 47742 20690
rect 47742 20638 47794 20690
rect 47794 20638 47796 20690
rect 47740 20636 47796 20638
rect 47628 19234 47684 19236
rect 47628 19182 47630 19234
rect 47630 19182 47682 19234
rect 47682 19182 47684 19234
rect 47628 19180 47684 19182
rect 46956 18956 47012 19012
rect 47068 18562 47124 18564
rect 47068 18510 47070 18562
rect 47070 18510 47122 18562
rect 47122 18510 47124 18562
rect 47068 18508 47124 18510
rect 47180 18450 47236 18452
rect 47180 18398 47182 18450
rect 47182 18398 47234 18450
rect 47234 18398 47236 18450
rect 47180 18396 47236 18398
rect 47068 17612 47124 17668
rect 46956 17442 47012 17444
rect 46956 17390 46958 17442
rect 46958 17390 47010 17442
rect 47010 17390 47012 17442
rect 46956 17388 47012 17390
rect 47628 17442 47684 17444
rect 47628 17390 47630 17442
rect 47630 17390 47682 17442
rect 47682 17390 47684 17442
rect 47628 17388 47684 17390
rect 47068 17106 47124 17108
rect 47068 17054 47070 17106
rect 47070 17054 47122 17106
rect 47122 17054 47124 17106
rect 47068 17052 47124 17054
rect 46732 15820 46788 15876
rect 47180 16044 47236 16100
rect 47068 15820 47124 15876
rect 46508 14812 46564 14868
rect 44940 10556 44996 10612
rect 45164 11452 45220 11508
rect 45164 10444 45220 10500
rect 45724 11452 45780 11508
rect 45052 10332 45108 10388
rect 44604 9996 44660 10052
rect 45276 9212 45332 9268
rect 44604 8876 44660 8932
rect 43932 8818 43988 8820
rect 43932 8766 43934 8818
rect 43934 8766 43986 8818
rect 43986 8766 43988 8818
rect 43932 8764 43988 8766
rect 43708 8428 43764 8484
rect 42476 7196 42532 7252
rect 44268 7420 44324 7476
rect 44940 8876 44996 8932
rect 45276 8428 45332 8484
rect 46508 14306 46564 14308
rect 46508 14254 46510 14306
rect 46510 14254 46562 14306
rect 46562 14254 46564 14306
rect 46508 14252 46564 14254
rect 46284 14140 46340 14196
rect 46060 13858 46116 13860
rect 46060 13806 46062 13858
rect 46062 13806 46114 13858
rect 46114 13806 46116 13858
rect 46060 13804 46116 13806
rect 46172 12290 46228 12292
rect 46172 12238 46174 12290
rect 46174 12238 46226 12290
rect 46226 12238 46228 12290
rect 46172 12236 46228 12238
rect 45836 10332 45892 10388
rect 46732 14418 46788 14420
rect 46732 14366 46734 14418
rect 46734 14366 46786 14418
rect 46786 14366 46788 14418
rect 46732 14364 46788 14366
rect 48972 18450 49028 18452
rect 48972 18398 48974 18450
rect 48974 18398 49026 18450
rect 49026 18398 49028 18450
rect 48972 18396 49028 18398
rect 49420 20524 49476 20580
rect 50540 21756 50596 21812
rect 50540 20914 50596 20916
rect 50540 20862 50542 20914
rect 50542 20862 50594 20914
rect 50594 20862 50596 20914
rect 50540 20860 50596 20862
rect 52892 22652 52948 22708
rect 53116 22316 53172 22372
rect 53228 22204 53284 22260
rect 57932 26236 57988 26292
rect 57932 24892 57988 24948
rect 55356 24220 55412 24276
rect 55580 23938 55636 23940
rect 55580 23886 55582 23938
rect 55582 23886 55634 23938
rect 55634 23886 55636 23938
rect 55580 23884 55636 23886
rect 54460 22316 54516 22372
rect 51548 21308 51604 21364
rect 51212 20860 51268 20916
rect 50540 20578 50596 20580
rect 50540 20526 50542 20578
rect 50542 20526 50594 20578
rect 50594 20526 50596 20578
rect 50540 20524 50596 20526
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 49644 20076 49700 20132
rect 49532 18396 49588 18452
rect 50540 19010 50596 19012
rect 50540 18958 50542 19010
rect 50542 18958 50594 19010
rect 50594 18958 50596 19010
rect 50540 18956 50596 18958
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 51100 18450 51156 18452
rect 51100 18398 51102 18450
rect 51102 18398 51154 18450
rect 51154 18398 51156 18450
rect 51100 18396 51156 18398
rect 51772 20914 51828 20916
rect 51772 20862 51774 20914
rect 51774 20862 51826 20914
rect 51826 20862 51828 20914
rect 51772 20860 51828 20862
rect 54236 22258 54292 22260
rect 54236 22206 54238 22258
rect 54238 22206 54290 22258
rect 54290 22206 54292 22258
rect 54236 22204 54292 22206
rect 53564 21420 53620 21476
rect 53340 20860 53396 20916
rect 54460 21474 54516 21476
rect 54460 21422 54462 21474
rect 54462 21422 54514 21474
rect 54514 21422 54516 21474
rect 54460 21420 54516 21422
rect 57932 20914 57988 20916
rect 57932 20862 57934 20914
rect 57934 20862 57986 20914
rect 57986 20862 57988 20914
rect 57932 20860 57988 20862
rect 51884 19180 51940 19236
rect 53228 19234 53284 19236
rect 53228 19182 53230 19234
rect 53230 19182 53282 19234
rect 53282 19182 53284 19234
rect 53228 19180 53284 19182
rect 52892 18956 52948 19012
rect 51660 18396 51716 18452
rect 47516 16098 47572 16100
rect 47516 16046 47518 16098
rect 47518 16046 47570 16098
rect 47570 16046 47572 16098
rect 47516 16044 47572 16046
rect 47964 17388 48020 17444
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 47964 17052 48020 17108
rect 48188 16604 48244 16660
rect 49532 16210 49588 16212
rect 49532 16158 49534 16210
rect 49534 16158 49586 16210
rect 49586 16158 49588 16210
rect 49532 16156 49588 16158
rect 50092 16156 50148 16212
rect 48076 15874 48132 15876
rect 48076 15822 48078 15874
rect 48078 15822 48130 15874
rect 48130 15822 48132 15874
rect 48076 15820 48132 15822
rect 49084 15820 49140 15876
rect 49644 15874 49700 15876
rect 49644 15822 49646 15874
rect 49646 15822 49698 15874
rect 49698 15822 49700 15874
rect 49644 15820 49700 15822
rect 48860 15036 48916 15092
rect 49420 15314 49476 15316
rect 49420 15262 49422 15314
rect 49422 15262 49474 15314
rect 49474 15262 49476 15314
rect 49420 15260 49476 15262
rect 49084 15148 49140 15204
rect 49980 15202 50036 15204
rect 49980 15150 49982 15202
rect 49982 15150 50034 15202
rect 50034 15150 50036 15202
rect 49980 15148 50036 15150
rect 49756 15036 49812 15092
rect 47180 13804 47236 13860
rect 46396 11506 46452 11508
rect 46396 11454 46398 11506
rect 46398 11454 46450 11506
rect 46450 11454 46452 11506
rect 46396 11452 46452 11454
rect 47404 12572 47460 12628
rect 46732 10668 46788 10724
rect 45612 9266 45668 9268
rect 45612 9214 45614 9266
rect 45614 9214 45666 9266
rect 45666 9214 45668 9266
rect 45612 9212 45668 9214
rect 48188 12124 48244 12180
rect 47516 11788 47572 11844
rect 46956 11394 47012 11396
rect 46956 11342 46958 11394
rect 46958 11342 47010 11394
rect 47010 11342 47012 11394
rect 46956 11340 47012 11342
rect 47292 10556 47348 10612
rect 50988 16156 51044 16212
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 51548 16828 51604 16884
rect 52668 18396 52724 18452
rect 53228 18508 53284 18564
rect 52108 17052 52164 17108
rect 53564 18396 53620 18452
rect 55132 18562 55188 18564
rect 55132 18510 55134 18562
rect 55134 18510 55186 18562
rect 55186 18510 55188 18562
rect 55132 18508 55188 18510
rect 54460 17106 54516 17108
rect 54460 17054 54462 17106
rect 54462 17054 54514 17106
rect 54514 17054 54516 17106
rect 54460 17052 54516 17054
rect 53340 16828 53396 16884
rect 52780 16604 52836 16660
rect 51772 16210 51828 16212
rect 51772 16158 51774 16210
rect 51774 16158 51826 16210
rect 51826 16158 51828 16210
rect 51772 16156 51828 16158
rect 51548 16098 51604 16100
rect 51548 16046 51550 16098
rect 51550 16046 51602 16098
rect 51602 16046 51604 16098
rect 51548 16044 51604 16046
rect 51212 15820 51268 15876
rect 53004 16210 53060 16212
rect 53004 16158 53006 16210
rect 53006 16158 53058 16210
rect 53058 16158 53060 16210
rect 53004 16156 53060 16158
rect 54572 16828 54628 16884
rect 54236 16658 54292 16660
rect 54236 16606 54238 16658
rect 54238 16606 54290 16658
rect 54290 16606 54292 16658
rect 54236 16604 54292 16606
rect 52892 16098 52948 16100
rect 52892 16046 52894 16098
rect 52894 16046 52946 16098
rect 52946 16046 52948 16098
rect 52892 16044 52948 16046
rect 52668 15426 52724 15428
rect 52668 15374 52670 15426
rect 52670 15374 52722 15426
rect 52722 15374 52724 15426
rect 52668 15372 52724 15374
rect 53564 15372 53620 15428
rect 50988 15314 51044 15316
rect 50988 15262 50990 15314
rect 50990 15262 51042 15314
rect 51042 15262 51044 15314
rect 50988 15260 51044 15262
rect 50876 14418 50932 14420
rect 50876 14366 50878 14418
rect 50878 14366 50930 14418
rect 50930 14366 50932 14418
rect 50876 14364 50932 14366
rect 51660 14364 51716 14420
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 52220 14364 52276 14420
rect 51660 13020 51716 13076
rect 51324 12962 51380 12964
rect 51324 12910 51326 12962
rect 51326 12910 51378 12962
rect 51378 12910 51380 12962
rect 51324 12908 51380 12910
rect 49756 12850 49812 12852
rect 49756 12798 49758 12850
rect 49758 12798 49810 12850
rect 49810 12798 49812 12850
rect 49756 12796 49812 12798
rect 48748 12348 48804 12404
rect 48972 12236 49028 12292
rect 48860 12178 48916 12180
rect 48860 12126 48862 12178
rect 48862 12126 48914 12178
rect 48914 12126 48916 12178
rect 48860 12124 48916 12126
rect 47628 11394 47684 11396
rect 47628 11342 47630 11394
rect 47630 11342 47682 11394
rect 47682 11342 47684 11394
rect 47628 11340 47684 11342
rect 46620 9826 46676 9828
rect 46620 9774 46622 9826
rect 46622 9774 46674 9826
rect 46674 9774 46676 9826
rect 46620 9772 46676 9774
rect 47964 10668 48020 10724
rect 48412 11788 48468 11844
rect 49308 12290 49364 12292
rect 49308 12238 49310 12290
rect 49310 12238 49362 12290
rect 49362 12238 49364 12290
rect 49308 12236 49364 12238
rect 50988 12684 51044 12740
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50204 12348 50260 12404
rect 49980 12290 50036 12292
rect 49980 12238 49982 12290
rect 49982 12238 50034 12290
rect 50034 12238 50036 12290
rect 49980 12236 50036 12238
rect 49532 12124 49588 12180
rect 49308 11394 49364 11396
rect 49308 11342 49310 11394
rect 49310 11342 49362 11394
rect 49362 11342 49364 11394
rect 49308 11340 49364 11342
rect 48076 10610 48132 10612
rect 48076 10558 48078 10610
rect 48078 10558 48130 10610
rect 48130 10558 48132 10610
rect 48076 10556 48132 10558
rect 48636 10556 48692 10612
rect 49644 10610 49700 10612
rect 49644 10558 49646 10610
rect 49646 10558 49698 10610
rect 49698 10558 49700 10610
rect 49644 10556 49700 10558
rect 50988 12236 51044 12292
rect 51100 12850 51156 12852
rect 51100 12798 51102 12850
rect 51102 12798 51154 12850
rect 51154 12798 51156 12850
rect 51100 12796 51156 12798
rect 51772 12796 51828 12852
rect 52780 13074 52836 13076
rect 52780 13022 52782 13074
rect 52782 13022 52834 13074
rect 52834 13022 52836 13074
rect 52780 13020 52836 13022
rect 53004 12962 53060 12964
rect 53004 12910 53006 12962
rect 53006 12910 53058 12962
rect 53058 12910 53060 12962
rect 53004 12908 53060 12910
rect 52108 12684 52164 12740
rect 51884 12402 51940 12404
rect 51884 12350 51886 12402
rect 51886 12350 51938 12402
rect 51938 12350 51940 12402
rect 51884 12348 51940 12350
rect 50764 12178 50820 12180
rect 50764 12126 50766 12178
rect 50766 12126 50818 12178
rect 50818 12126 50820 12178
rect 50764 12124 50820 12126
rect 52668 12348 52724 12404
rect 54572 14476 54628 14532
rect 55580 14530 55636 14532
rect 55580 14478 55582 14530
rect 55582 14478 55634 14530
rect 55634 14478 55636 14530
rect 55580 14476 55636 14478
rect 52332 12124 52388 12180
rect 52108 11676 52164 11732
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 53452 12178 53508 12180
rect 53452 12126 53454 12178
rect 53454 12126 53506 12178
rect 53506 12126 53508 12178
rect 53452 12124 53508 12126
rect 53900 12124 53956 12180
rect 52780 11676 52836 11732
rect 52220 11340 52276 11396
rect 50428 10556 50484 10612
rect 50092 10332 50148 10388
rect 46284 9212 46340 9268
rect 50540 10332 50596 10388
rect 51100 10610 51156 10612
rect 51100 10558 51102 10610
rect 51102 10558 51154 10610
rect 51154 10558 51156 10610
rect 51100 10556 51156 10558
rect 50764 10498 50820 10500
rect 50764 10446 50766 10498
rect 50766 10446 50818 10498
rect 50818 10446 50820 10498
rect 50764 10444 50820 10446
rect 51212 10332 51268 10388
rect 50204 9660 50260 9716
rect 51660 9714 51716 9716
rect 51660 9662 51662 9714
rect 51662 9662 51714 9714
rect 51714 9662 51716 9714
rect 51660 9660 51716 9662
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 47852 9100 47908 9156
rect 45500 8316 45556 8372
rect 47740 8316 47796 8372
rect 43932 7308 43988 7364
rect 45500 7474 45556 7476
rect 45500 7422 45502 7474
rect 45502 7422 45554 7474
rect 45554 7422 45556 7474
rect 45500 7420 45556 7422
rect 45276 7308 45332 7364
rect 43484 6690 43540 6692
rect 43484 6638 43486 6690
rect 43486 6638 43538 6690
rect 43538 6638 43540 6690
rect 43484 6636 43540 6638
rect 42140 5964 42196 6020
rect 46284 7420 46340 7476
rect 46172 7196 46228 7252
rect 48860 9154 48916 9156
rect 48860 9102 48862 9154
rect 48862 9102 48914 9154
rect 48914 9102 48916 9154
rect 48860 9100 48916 9102
rect 49308 8316 49364 8372
rect 48412 8034 48468 8036
rect 48412 7982 48414 8034
rect 48414 7982 48466 8034
rect 48466 7982 48468 8034
rect 48412 7980 48468 7982
rect 48972 7980 49028 8036
rect 49308 7474 49364 7476
rect 49308 7422 49310 7474
rect 49310 7422 49362 7474
rect 49362 7422 49364 7474
rect 49308 7420 49364 7422
rect 47964 7196 48020 7252
rect 46732 6524 46788 6580
rect 49196 7250 49252 7252
rect 49196 7198 49198 7250
rect 49198 7198 49250 7250
rect 49250 7198 49252 7250
rect 49196 7196 49252 7198
rect 51996 8988 52052 9044
rect 49532 8316 49588 8372
rect 51548 8876 51604 8932
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 53788 11676 53844 11732
rect 54572 12178 54628 12180
rect 54572 12126 54574 12178
rect 54574 12126 54626 12178
rect 54626 12126 54628 12178
rect 54572 12124 54628 12126
rect 54348 11788 54404 11844
rect 57932 17500 57988 17556
rect 57932 14812 57988 14868
rect 57932 12124 57988 12180
rect 55692 11788 55748 11844
rect 54236 11394 54292 11396
rect 54236 11342 54238 11394
rect 54238 11342 54290 11394
rect 54290 11342 54292 11394
rect 54236 11340 54292 11342
rect 52668 9042 52724 9044
rect 52668 8990 52670 9042
rect 52670 8990 52722 9042
rect 52722 8990 52724 9042
rect 52668 8988 52724 8990
rect 52556 8930 52612 8932
rect 52556 8878 52558 8930
rect 52558 8878 52610 8930
rect 52610 8878 52612 8930
rect 52556 8876 52612 8878
rect 57932 8370 57988 8372
rect 57932 8318 57934 8370
rect 57934 8318 57986 8370
rect 57986 8318 57988 8370
rect 57932 8316 57988 8318
rect 54012 8204 54068 8260
rect 55580 8258 55636 8260
rect 55580 8206 55582 8258
rect 55582 8206 55634 8258
rect 55634 8206 55636 8258
rect 55580 8204 55636 8206
rect 49868 6748 49924 6804
rect 50540 6802 50596 6804
rect 50540 6750 50542 6802
rect 50542 6750 50594 6802
rect 50594 6750 50596 6802
rect 50540 6748 50596 6750
rect 51436 7474 51492 7476
rect 51436 7422 51438 7474
rect 51438 7422 51490 7474
rect 51490 7422 51492 7474
rect 51436 7420 51492 7422
rect 50652 6690 50708 6692
rect 50652 6638 50654 6690
rect 50654 6638 50706 6690
rect 50706 6638 50708 6690
rect 50652 6636 50708 6638
rect 47964 6300 48020 6356
rect 46508 6018 46564 6020
rect 46508 5966 46510 6018
rect 46510 5966 46562 6018
rect 46562 5966 46564 6018
rect 46508 5964 46564 5966
rect 42588 5068 42644 5124
rect 42812 5180 42868 5236
rect 45388 5180 45444 5236
rect 43372 5122 43428 5124
rect 43372 5070 43374 5122
rect 43374 5070 43426 5122
rect 43426 5070 43428 5122
rect 43372 5068 43428 5070
rect 45164 5122 45220 5124
rect 45164 5070 45166 5122
rect 45166 5070 45218 5122
rect 45218 5070 45220 5122
rect 45164 5068 45220 5070
rect 41244 5010 41300 5012
rect 41244 4958 41246 5010
rect 41246 4958 41298 5010
rect 41298 4958 41300 5010
rect 41244 4956 41300 4958
rect 46172 5180 46228 5236
rect 40348 4338 40404 4340
rect 40348 4286 40350 4338
rect 40350 4286 40402 4338
rect 40402 4286 40404 4338
rect 40348 4284 40404 4286
rect 41132 4338 41188 4340
rect 41132 4286 41134 4338
rect 41134 4286 41186 4338
rect 41186 4286 41188 4338
rect 41132 4284 41188 4286
rect 46396 5068 46452 5124
rect 47180 6018 47236 6020
rect 47180 5966 47182 6018
rect 47182 5966 47234 6018
rect 47234 5966 47236 6018
rect 47180 5964 47236 5966
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 43708 3388 43764 3444
rect 39116 3164 39172 3220
rect 39004 1484 39060 1540
rect 7868 1372 7924 1428
rect 44940 3388 44996 3444
rect 51772 3612 51828 3668
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 58156 5404 58212 5460
rect 58156 4732 58212 4788
rect 58156 4060 58212 4116
rect 52892 3666 52948 3668
rect 52892 3614 52894 3666
rect 52894 3614 52946 3666
rect 52946 3614 52948 3666
rect 52892 3612 52948 3614
rect 58156 3330 58212 3332
rect 58156 3278 58158 3330
rect 58158 3278 58210 3330
rect 58210 3278 58212 3330
rect 58156 3276 58212 3278
rect 57708 2716 57764 2772
<< metal3 >>
rect 15362 57148 15372 57204
rect 15428 57148 28140 57204
rect 28196 57148 28206 57204
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 47730 56252 47740 56308
rect 47796 56252 48972 56308
rect 49028 56252 49038 56308
rect 49186 56252 49196 56308
rect 49252 56252 52220 56308
rect 52276 56252 52286 56308
rect 53106 56252 53116 56308
rect 53172 56252 54124 56308
rect 54180 56252 54190 56308
rect 54450 56252 54460 56308
rect 54516 56252 55468 56308
rect 55524 56252 55534 56308
rect 30370 56028 30380 56084
rect 30436 56028 31164 56084
rect 31220 56028 32284 56084
rect 32340 56028 32350 56084
rect 49522 56028 49532 56084
rect 49588 56028 51212 56084
rect 51268 56028 51278 56084
rect 33506 55916 33516 55972
rect 33572 55916 34860 55972
rect 34916 55916 34926 55972
rect 55122 55916 55132 55972
rect 55188 55916 55916 55972
rect 55972 55916 55982 55972
rect 59200 55860 60000 55888
rect 58146 55804 58156 55860
rect 58212 55804 60000 55860
rect 59200 55776 60000 55804
rect 18050 55692 18060 55748
rect 18116 55692 31612 55748
rect 31668 55692 31678 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 15810 55580 15820 55636
rect 15876 55580 28588 55636
rect 28644 55580 28654 55636
rect 20962 55468 20972 55524
rect 21028 55468 28700 55524
rect 28756 55468 28766 55524
rect 48402 55356 48412 55412
rect 48468 55356 49644 55412
rect 49700 55356 49710 55412
rect 52434 55356 52444 55412
rect 52500 55356 53676 55412
rect 53732 55356 53742 55412
rect 31892 55244 33068 55300
rect 33124 55244 33134 55300
rect 34066 55244 34076 55300
rect 34132 55244 36988 55300
rect 37044 55244 37054 55300
rect 31892 55188 31948 55244
rect 59200 55188 60000 55216
rect 19180 55132 19964 55188
rect 20020 55132 20030 55188
rect 30146 55132 30156 55188
rect 30212 55132 30828 55188
rect 30884 55132 30894 55188
rect 31490 55132 31500 55188
rect 31556 55132 31948 55188
rect 33842 55132 33852 55188
rect 33908 55132 33918 55188
rect 41010 55132 41020 55188
rect 41076 55132 42476 55188
rect 42532 55132 42542 55188
rect 42914 55132 42924 55188
rect 42980 55132 44828 55188
rect 44884 55132 45500 55188
rect 45556 55132 45566 55188
rect 45714 55132 45724 55188
rect 45780 55132 47068 55188
rect 47124 55132 47134 55188
rect 57698 55132 57708 55188
rect 57764 55132 60000 55188
rect 19180 55076 19236 55132
rect 18722 55020 18732 55076
rect 18788 55020 19180 55076
rect 19236 55020 19246 55076
rect 19842 55020 19852 55076
rect 19908 55020 23324 55076
rect 23380 55020 23390 55076
rect 27430 55020 27468 55076
rect 27524 55020 27534 55076
rect 27906 55020 27916 55076
rect 27972 55020 30604 55076
rect 30660 55020 30670 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 22194 54796 22204 54852
rect 22260 54796 22764 54852
rect 22820 54796 22830 54852
rect 24882 54796 24892 54852
rect 24948 54796 28588 54852
rect 28644 54796 29372 54852
rect 29428 54796 29438 54852
rect 33852 54740 33908 55132
rect 59200 55104 60000 55132
rect 42130 55020 42140 55076
rect 42196 55020 44940 55076
rect 44996 55020 45006 55076
rect 45154 55020 45164 55076
rect 45220 55020 49084 55076
rect 49140 55020 49980 55076
rect 50036 55020 50046 55076
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 51090 54796 51100 54852
rect 51156 54796 52332 54852
rect 52388 54796 52398 54852
rect 17826 54684 17836 54740
rect 17892 54684 28028 54740
rect 28084 54684 28094 54740
rect 33842 54684 33852 54740
rect 33908 54684 33918 54740
rect 21634 54572 21644 54628
rect 21700 54572 22428 54628
rect 22484 54572 23660 54628
rect 23716 54572 23726 54628
rect 29474 54572 29484 54628
rect 29540 54572 31948 54628
rect 32004 54572 33180 54628
rect 33236 54572 33246 54628
rect 46834 54572 46844 54628
rect 46900 54572 47628 54628
rect 47684 54572 47694 54628
rect 59200 54516 60000 54544
rect 20402 54460 20412 54516
rect 20468 54460 21420 54516
rect 21476 54460 22204 54516
rect 22260 54460 22270 54516
rect 23314 54460 23324 54516
rect 23380 54460 25116 54516
rect 25172 54460 25182 54516
rect 25890 54460 25900 54516
rect 25956 54460 27132 54516
rect 27188 54460 29708 54516
rect 29764 54460 29774 54516
rect 42242 54460 42252 54516
rect 42308 54460 43484 54516
rect 43540 54460 43550 54516
rect 44370 54460 44380 54516
rect 44436 54460 49308 54516
rect 49364 54460 50092 54516
rect 50148 54460 50158 54516
rect 58146 54460 58156 54516
rect 58212 54460 60000 54516
rect 59200 54432 60000 54460
rect 19058 54348 19068 54404
rect 19124 54348 21196 54404
rect 21252 54348 21262 54404
rect 21522 54348 21532 54404
rect 21588 54348 25676 54404
rect 25732 54348 25742 54404
rect 30146 54348 30156 54404
rect 30212 54348 34076 54404
rect 34132 54348 35420 54404
rect 35476 54348 35486 54404
rect 37762 54348 37772 54404
rect 37828 54348 38444 54404
rect 38500 54348 39900 54404
rect 39956 54348 39966 54404
rect 19842 54236 19852 54292
rect 19908 54236 21308 54292
rect 21364 54236 25564 54292
rect 25620 54236 25630 54292
rect 27234 54236 27244 54292
rect 27300 54236 33852 54292
rect 33908 54236 33918 54292
rect 35186 54236 35196 54292
rect 35252 54236 42588 54292
rect 42644 54236 42654 54292
rect 20860 54124 22652 54180
rect 22708 54124 22718 54180
rect 22866 54124 22876 54180
rect 22932 54124 26908 54180
rect 46946 54124 46956 54180
rect 47012 54124 47516 54180
rect 47572 54124 50876 54180
rect 50932 54124 50942 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 20860 54068 20916 54124
rect 26852 54068 26908 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 19516 54012 20860 54068
rect 20916 54012 20926 54068
rect 26852 54012 27804 54068
rect 27860 54012 27870 54068
rect 0 53844 800 53872
rect 19516 53844 19572 54012
rect 19740 53900 24164 53956
rect 25554 53900 25564 53956
rect 25620 53900 30044 53956
rect 30100 53900 30110 53956
rect 39778 53900 39788 53956
rect 39844 53900 46172 53956
rect 46228 53900 46238 53956
rect 19740 53844 19796 53900
rect 0 53788 1708 53844
rect 1764 53788 1774 53844
rect 16930 53788 16940 53844
rect 16996 53788 17836 53844
rect 17892 53788 17902 53844
rect 19506 53788 19516 53844
rect 19572 53788 19582 53844
rect 19730 53788 19740 53844
rect 19796 53788 19806 53844
rect 22306 53788 22316 53844
rect 22372 53788 23884 53844
rect 23940 53788 23950 53844
rect 0 53760 800 53788
rect 24108 53732 24164 53900
rect 25218 53788 25228 53844
rect 25284 53788 25788 53844
rect 25844 53788 25854 53844
rect 28466 53788 28476 53844
rect 28532 53788 30940 53844
rect 30996 53788 31006 53844
rect 37986 53788 37996 53844
rect 38052 53788 41356 53844
rect 41412 53788 41422 53844
rect 43586 53788 43596 53844
rect 43652 53788 43820 53844
rect 43876 53788 43886 53844
rect 19618 53676 19628 53732
rect 19684 53676 20300 53732
rect 20356 53676 20366 53732
rect 22530 53676 22540 53732
rect 22596 53676 23436 53732
rect 23492 53676 23502 53732
rect 24108 53676 31948 53732
rect 32004 53676 32014 53732
rect 34402 53676 34412 53732
rect 34468 53676 36092 53732
rect 36148 53676 37324 53732
rect 37380 53676 37390 53732
rect 47170 53676 47180 53732
rect 47236 53676 47852 53732
rect 47908 53676 47918 53732
rect 50082 53676 50092 53732
rect 50148 53676 50988 53732
rect 51044 53676 51054 53732
rect 16034 53564 16044 53620
rect 16100 53564 16716 53620
rect 16772 53564 16782 53620
rect 33282 53564 33292 53620
rect 33348 53564 35084 53620
rect 35140 53564 35150 53620
rect 35858 53564 35868 53620
rect 35924 53564 37212 53620
rect 37268 53564 37278 53620
rect 38098 53564 38108 53620
rect 38164 53564 39452 53620
rect 39508 53564 39518 53620
rect 43922 53564 43932 53620
rect 43988 53564 44828 53620
rect 44884 53564 49644 53620
rect 49700 53564 49710 53620
rect 51650 53564 51660 53620
rect 51716 53564 52668 53620
rect 52724 53564 52734 53620
rect 14914 53452 14924 53508
rect 14980 53452 16492 53508
rect 16548 53452 17500 53508
rect 17556 53452 20412 53508
rect 20468 53452 20478 53508
rect 20710 53452 20748 53508
rect 20804 53452 22316 53508
rect 22372 53452 23324 53508
rect 23380 53452 23390 53508
rect 25890 53452 25900 53508
rect 25956 53452 26908 53508
rect 26964 53452 26974 53508
rect 27682 53452 27692 53508
rect 27748 53452 28252 53508
rect 28308 53452 28318 53508
rect 36418 53452 36428 53508
rect 36484 53452 42028 53508
rect 42084 53452 42094 53508
rect 50306 53452 50316 53508
rect 50372 53452 51324 53508
rect 51380 53452 51390 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 17154 53228 17164 53284
rect 17220 53228 18844 53284
rect 18900 53228 18910 53284
rect 19394 53228 19404 53284
rect 19460 53228 19628 53284
rect 19684 53228 19694 53284
rect 20514 53228 20524 53284
rect 20580 53228 23436 53284
rect 23492 53228 25340 53284
rect 25396 53228 25406 53284
rect 26786 53228 26796 53284
rect 26852 53228 28140 53284
rect 28196 53228 28812 53284
rect 28868 53228 28878 53284
rect 20524 53172 20580 53228
rect 17714 53116 17724 53172
rect 17780 53116 18900 53172
rect 19282 53116 19292 53172
rect 19348 53116 20580 53172
rect 22754 53116 22764 53172
rect 22820 53116 23100 53172
rect 23156 53116 23166 53172
rect 25106 53116 25116 53172
rect 25172 53116 30828 53172
rect 30884 53116 30894 53172
rect 18844 53060 18900 53116
rect 17490 53004 17500 53060
rect 17556 53004 18620 53060
rect 18676 53004 18686 53060
rect 18844 53004 28588 53060
rect 28644 53004 28654 53060
rect 49186 53004 49196 53060
rect 49252 53004 50652 53060
rect 50708 53004 50718 53060
rect 17602 52892 17612 52948
rect 17668 52892 19068 52948
rect 19124 52892 19134 52948
rect 19628 52892 21756 52948
rect 21812 52892 21822 52948
rect 21970 52892 21980 52948
rect 22036 52892 22540 52948
rect 22596 52892 22606 52948
rect 23202 52892 23212 52948
rect 23268 52892 32116 52948
rect 32946 52892 32956 52948
rect 33012 52892 34300 52948
rect 34356 52892 34748 52948
rect 34804 52892 34814 52948
rect 34962 52892 34972 52948
rect 35028 52892 36316 52948
rect 36372 52892 37100 52948
rect 37156 52892 37166 52948
rect 19628 52836 19684 52892
rect 18386 52780 18396 52836
rect 18452 52780 19684 52836
rect 19842 52780 19852 52836
rect 19908 52780 21196 52836
rect 21252 52780 21262 52836
rect 30930 52780 30940 52836
rect 30996 52780 31948 52836
rect 15586 52668 15596 52724
rect 15652 52668 26908 52724
rect 30370 52668 30380 52724
rect 30436 52668 31164 52724
rect 31220 52668 31724 52724
rect 31780 52668 31790 52724
rect 26852 52612 26908 52668
rect 16930 52556 16940 52612
rect 16996 52556 18172 52612
rect 18228 52556 18238 52612
rect 19170 52556 19180 52612
rect 19236 52556 19964 52612
rect 20020 52556 20030 52612
rect 26852 52556 30156 52612
rect 30212 52556 30222 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 20300 52444 20524 52500
rect 20580 52444 21196 52500
rect 21252 52444 21262 52500
rect 21420 52444 25564 52500
rect 25620 52444 26460 52500
rect 26516 52444 26908 52500
rect 20300 52276 20356 52444
rect 21420 52388 21476 52444
rect 20626 52332 20636 52388
rect 20692 52332 21420 52388
rect 21476 52332 21486 52388
rect 22978 52332 22988 52388
rect 23044 52332 23212 52388
rect 23268 52332 23278 52388
rect 26852 52276 26908 52444
rect 14130 52220 14140 52276
rect 14196 52220 18284 52276
rect 18340 52220 18350 52276
rect 19394 52220 19404 52276
rect 19460 52220 20356 52276
rect 21298 52220 21308 52276
rect 21364 52220 22092 52276
rect 22148 52220 22158 52276
rect 23090 52220 23100 52276
rect 23156 52220 25340 52276
rect 25396 52220 25406 52276
rect 26852 52220 27356 52276
rect 27412 52220 27422 52276
rect 18050 52108 18060 52164
rect 18116 52108 19180 52164
rect 19236 52108 19246 52164
rect 20850 52108 20860 52164
rect 20916 52108 21868 52164
rect 21924 52108 21934 52164
rect 23986 52108 23996 52164
rect 24052 52108 26908 52164
rect 26964 52108 26974 52164
rect 31892 52052 31948 52780
rect 32060 52724 32116 52892
rect 32274 52780 32284 52836
rect 32340 52780 34076 52836
rect 34132 52780 34636 52836
rect 34692 52780 34702 52836
rect 32060 52668 38444 52724
rect 38500 52668 38510 52724
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 59200 52500 60000 52528
rect 58146 52444 58156 52500
rect 58212 52444 60000 52500
rect 59200 52416 60000 52444
rect 34850 52332 34860 52388
rect 34916 52332 38108 52388
rect 38164 52332 38174 52388
rect 35074 52108 35084 52164
rect 35140 52108 42252 52164
rect 42308 52108 42318 52164
rect 42578 52108 42588 52164
rect 42644 52108 43932 52164
rect 43988 52108 44940 52164
rect 44996 52108 45006 52164
rect 51426 52108 51436 52164
rect 51492 52108 51502 52164
rect 51436 52052 51492 52108
rect 17154 51996 17164 52052
rect 17220 51996 20524 52052
rect 20580 51996 20590 52052
rect 22306 51996 22316 52052
rect 22372 51996 23772 52052
rect 23828 51996 23838 52052
rect 25330 51996 25340 52052
rect 25396 51996 27692 52052
rect 27748 51996 27758 52052
rect 30818 51996 30828 52052
rect 30884 51996 31276 52052
rect 31332 51996 31342 52052
rect 31892 51996 38780 52052
rect 38836 51996 38846 52052
rect 51090 51996 51100 52052
rect 51156 51996 51492 52052
rect 23874 51884 23884 51940
rect 23940 51884 25004 51940
rect 25060 51884 25070 51940
rect 27234 51884 27244 51940
rect 27300 51884 37548 51940
rect 37604 51884 37614 51940
rect 39442 51884 39452 51940
rect 39508 51884 40796 51940
rect 40852 51884 40862 51940
rect 19590 51772 19628 51828
rect 19684 51772 19694 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 22988 51660 31164 51716
rect 31220 51660 31230 51716
rect 41010 51660 41020 51716
rect 41076 51660 42140 51716
rect 42196 51660 43148 51716
rect 43204 51660 43214 51716
rect 22988 51604 23044 51660
rect 15474 51548 15484 51604
rect 15540 51548 16716 51604
rect 16772 51548 16782 51604
rect 22978 51548 22988 51604
rect 23044 51548 23054 51604
rect 23874 51548 23884 51604
rect 23940 51548 24892 51604
rect 24948 51548 24958 51604
rect 25666 51548 25676 51604
rect 25732 51548 31948 51604
rect 23622 51436 23660 51492
rect 23716 51436 23726 51492
rect 24994 51436 25004 51492
rect 25060 51436 28252 51492
rect 28308 51436 29260 51492
rect 29316 51436 29326 51492
rect 30930 51436 30940 51492
rect 30996 51436 31164 51492
rect 31220 51436 31230 51492
rect 31892 51380 31948 51548
rect 36978 51436 36988 51492
rect 37044 51436 42028 51492
rect 42084 51436 42094 51492
rect 46050 51436 46060 51492
rect 46116 51436 46844 51492
rect 46900 51436 47404 51492
rect 47460 51436 47470 51492
rect 16258 51324 16268 51380
rect 16324 51324 17556 51380
rect 18386 51324 18396 51380
rect 18452 51324 18844 51380
rect 18900 51324 18910 51380
rect 19170 51324 19180 51380
rect 19236 51324 22484 51380
rect 22642 51324 22652 51380
rect 22708 51324 24108 51380
rect 24164 51324 24174 51380
rect 25330 51324 25340 51380
rect 25396 51324 25788 51380
rect 25844 51324 25854 51380
rect 26450 51324 26460 51380
rect 26516 51324 28364 51380
rect 28420 51324 28430 51380
rect 30146 51324 30156 51380
rect 30212 51324 30828 51380
rect 30884 51324 30894 51380
rect 31892 51324 36092 51380
rect 36148 51324 36158 51380
rect 38546 51324 38556 51380
rect 38612 51324 39116 51380
rect 39172 51324 39182 51380
rect 40002 51324 40012 51380
rect 40068 51324 41132 51380
rect 41188 51324 41198 51380
rect 51202 51324 51212 51380
rect 51268 51324 52332 51380
rect 52388 51324 52398 51380
rect 17500 51268 17556 51324
rect 22428 51268 22484 51324
rect 15474 51212 15484 51268
rect 15540 51212 16380 51268
rect 16436 51212 16446 51268
rect 17490 51212 17500 51268
rect 17556 51212 18284 51268
rect 18340 51212 18350 51268
rect 19282 51212 19292 51268
rect 19348 51212 21756 51268
rect 21812 51212 21822 51268
rect 22428 51212 22988 51268
rect 23044 51212 23054 51268
rect 24994 51212 25004 51268
rect 25060 51212 30716 51268
rect 30772 51212 30782 51268
rect 31154 51212 31164 51268
rect 31220 51212 34076 51268
rect 34132 51212 34142 51268
rect 44034 51212 44044 51268
rect 44100 51212 50428 51268
rect 50484 51212 51548 51268
rect 51604 51212 51614 51268
rect 59200 51156 60000 51184
rect 11890 51100 11900 51156
rect 11956 51100 18396 51156
rect 18452 51100 20188 51156
rect 20244 51100 22540 51156
rect 22596 51100 22606 51156
rect 23874 51100 23884 51156
rect 23940 51100 25564 51156
rect 25620 51100 25630 51156
rect 25788 51100 27244 51156
rect 27300 51100 27310 51156
rect 31378 51100 31388 51156
rect 31444 51100 33180 51156
rect 33236 51100 33246 51156
rect 34738 51100 34748 51156
rect 34804 51100 37660 51156
rect 37716 51100 37726 51156
rect 37874 51100 37884 51156
rect 37940 51100 38780 51156
rect 38836 51100 38846 51156
rect 39218 51100 39228 51156
rect 39284 51100 40908 51156
rect 40964 51100 40974 51156
rect 57922 51100 57932 51156
rect 57988 51100 60000 51156
rect 25788 51044 25844 51100
rect 59200 51072 60000 51100
rect 14354 50988 14364 51044
rect 14420 50988 18732 51044
rect 18788 50988 18798 51044
rect 19618 50988 19628 51044
rect 19684 50988 23212 51044
rect 23268 50988 25844 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 15698 50876 15708 50932
rect 15764 50876 16604 50932
rect 16660 50876 25228 50932
rect 25284 50876 25294 50932
rect 44258 50876 44268 50932
rect 44324 50876 45500 50932
rect 45556 50876 45566 50932
rect 18386 50764 18396 50820
rect 18452 50764 19628 50820
rect 19684 50764 19694 50820
rect 20934 50764 20972 50820
rect 21028 50764 21038 50820
rect 12002 50652 12012 50708
rect 12068 50652 12908 50708
rect 12964 50652 13468 50708
rect 13524 50652 17388 50708
rect 17444 50652 17454 50708
rect 18946 50652 18956 50708
rect 19012 50652 19516 50708
rect 19572 50652 19582 50708
rect 22764 50652 26516 50708
rect 27570 50652 27580 50708
rect 27636 50652 28252 50708
rect 28308 50652 28318 50708
rect 38322 50652 38332 50708
rect 38388 50652 39004 50708
rect 39060 50652 39788 50708
rect 39844 50652 39854 50708
rect 15586 50540 15596 50596
rect 15652 50540 19012 50596
rect 14578 50428 14588 50484
rect 14644 50428 15260 50484
rect 15316 50428 15326 50484
rect 18956 50372 19012 50540
rect 19404 50540 22092 50596
rect 22148 50540 22158 50596
rect 22306 50540 22316 50596
rect 22372 50540 22410 50596
rect 19404 50372 19460 50540
rect 22764 50484 22820 50652
rect 23202 50540 23212 50596
rect 23268 50540 23996 50596
rect 24052 50540 24062 50596
rect 25526 50540 25564 50596
rect 25620 50540 25630 50596
rect 26460 50484 26516 50652
rect 27346 50540 27356 50596
rect 27412 50540 27804 50596
rect 27860 50540 27870 50596
rect 29138 50540 29148 50596
rect 29204 50540 30044 50596
rect 30100 50540 30110 50596
rect 33282 50540 33292 50596
rect 33348 50540 33964 50596
rect 34020 50540 34030 50596
rect 37538 50540 37548 50596
rect 37604 50540 39340 50596
rect 39396 50540 39406 50596
rect 42466 50540 42476 50596
rect 42532 50540 43036 50596
rect 43092 50540 43484 50596
rect 43540 50540 43550 50596
rect 47954 50540 47964 50596
rect 48020 50540 48636 50596
rect 48692 50540 48702 50596
rect 50978 50540 50988 50596
rect 51044 50540 51660 50596
rect 51716 50540 52892 50596
rect 52948 50540 52958 50596
rect 53890 50540 53900 50596
rect 53956 50540 55580 50596
rect 55636 50540 55646 50596
rect 20850 50428 20860 50484
rect 20916 50428 21868 50484
rect 21924 50428 21934 50484
rect 22642 50428 22652 50484
rect 22708 50428 22820 50484
rect 23090 50428 23100 50484
rect 23156 50428 23548 50484
rect 26450 50428 26460 50484
rect 26516 50428 26908 50484
rect 26964 50428 26974 50484
rect 28130 50428 28140 50484
rect 28196 50428 28476 50484
rect 28532 50428 28542 50484
rect 31826 50428 31836 50484
rect 31892 50428 32956 50484
rect 33012 50428 33022 50484
rect 38994 50428 39004 50484
rect 39060 50428 39900 50484
rect 39956 50428 39966 50484
rect 44146 50428 44156 50484
rect 44212 50428 45164 50484
rect 45220 50428 45230 50484
rect 45388 50428 46620 50484
rect 46676 50428 47068 50484
rect 47124 50428 47134 50484
rect 50642 50428 50652 50484
rect 50708 50428 51100 50484
rect 51156 50428 51166 50484
rect 51874 50428 51884 50484
rect 51940 50428 52780 50484
rect 52836 50428 52846 50484
rect 58146 50428 58156 50484
rect 58212 50428 59332 50484
rect 23492 50372 23548 50428
rect 44156 50372 44212 50428
rect 45388 50372 45444 50428
rect 15138 50316 15148 50372
rect 15204 50316 15708 50372
rect 15764 50316 15774 50372
rect 18956 50316 19460 50372
rect 20290 50316 20300 50372
rect 20356 50316 21420 50372
rect 21476 50316 21486 50372
rect 23492 50316 27356 50372
rect 27412 50316 27422 50372
rect 28802 50316 28812 50372
rect 28868 50316 29708 50372
rect 29764 50316 30268 50372
rect 30324 50316 30334 50372
rect 30454 50316 30492 50372
rect 30548 50316 30558 50372
rect 31042 50316 31052 50372
rect 31108 50316 31500 50372
rect 31556 50316 31566 50372
rect 38612 50316 44212 50372
rect 44482 50316 44492 50372
rect 44548 50316 45444 50372
rect 38612 50260 38668 50316
rect 15474 50204 15484 50260
rect 15540 50204 19516 50260
rect 19572 50204 19582 50260
rect 36866 50204 36876 50260
rect 36932 50204 38668 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 16706 50092 16716 50148
rect 16772 50092 17052 50148
rect 17108 50092 17118 50148
rect 18918 50092 18956 50148
rect 19012 50092 19022 50148
rect 59276 50036 59332 50428
rect 18610 49980 18620 50036
rect 18676 49980 19404 50036
rect 19460 49980 19470 50036
rect 21074 49980 21084 50036
rect 21140 49980 35420 50036
rect 35476 49980 38108 50036
rect 38164 49980 38174 50036
rect 59052 49980 59332 50036
rect 12460 49868 17836 49924
rect 17892 49868 17902 49924
rect 18610 49868 18620 49924
rect 18676 49868 19628 49924
rect 19684 49868 23996 49924
rect 24052 49868 24062 49924
rect 27122 49868 27132 49924
rect 27188 49868 30044 49924
rect 30100 49868 30110 49924
rect 37650 49868 37660 49924
rect 37716 49868 43036 49924
rect 43092 49868 43102 49924
rect 12460 49700 12516 49868
rect 59052 49812 59108 49980
rect 59200 49812 60000 49840
rect 15250 49756 15260 49812
rect 15316 49756 16380 49812
rect 16436 49756 17500 49812
rect 17556 49756 19236 49812
rect 21746 49756 21756 49812
rect 21812 49756 22428 49812
rect 22484 49756 22494 49812
rect 22642 49756 22652 49812
rect 22708 49756 24108 49812
rect 24164 49756 28028 49812
rect 28084 49756 28094 49812
rect 30258 49756 30268 49812
rect 30324 49756 30716 49812
rect 30772 49756 30782 49812
rect 35634 49756 35644 49812
rect 35700 49756 36428 49812
rect 36484 49756 36494 49812
rect 43362 49756 43372 49812
rect 43428 49756 49868 49812
rect 49924 49756 49934 49812
rect 59052 49756 60000 49812
rect 19180 49700 19236 49756
rect 59200 49728 60000 49756
rect 11666 49644 11676 49700
rect 11732 49644 12124 49700
rect 12180 49644 12292 49700
rect 12450 49644 12460 49700
rect 12516 49644 12526 49700
rect 13458 49644 13468 49700
rect 13524 49644 14700 49700
rect 14756 49644 14766 49700
rect 16818 49644 16828 49700
rect 16884 49644 18956 49700
rect 19012 49644 19022 49700
rect 19180 49644 24052 49700
rect 24210 49644 24220 49700
rect 24276 49644 25228 49700
rect 25284 49644 26684 49700
rect 26740 49644 26750 49700
rect 26852 49644 27916 49700
rect 27972 49644 28588 49700
rect 28644 49644 29708 49700
rect 29764 49644 29774 49700
rect 35410 49644 35420 49700
rect 35476 49644 37436 49700
rect 37492 49644 37502 49700
rect 37986 49644 37996 49700
rect 38052 49644 50092 49700
rect 50148 49644 50158 49700
rect 11218 49532 11228 49588
rect 11284 49532 12012 49588
rect 12068 49532 12078 49588
rect 12236 49476 12292 49644
rect 23996 49588 24052 49644
rect 26852 49588 26908 49644
rect 14018 49532 14028 49588
rect 14084 49532 20188 49588
rect 20244 49532 20524 49588
rect 20580 49532 20590 49588
rect 21186 49532 21196 49588
rect 21252 49532 22428 49588
rect 22484 49532 22494 49588
rect 22978 49532 22988 49588
rect 23044 49532 23772 49588
rect 23828 49532 23838 49588
rect 23996 49532 26908 49588
rect 45378 49532 45388 49588
rect 45444 49532 46172 49588
rect 46228 49532 46238 49588
rect 12236 49420 14588 49476
rect 14644 49420 24668 49476
rect 24724 49420 25228 49476
rect 25284 49420 25294 49476
rect 26898 49420 26908 49476
rect 26964 49420 29148 49476
rect 29204 49420 29214 49476
rect 31042 49420 31052 49476
rect 31108 49420 31612 49476
rect 31668 49420 31678 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 14466 49308 14476 49364
rect 14532 49308 16940 49364
rect 16996 49308 17836 49364
rect 17892 49308 29260 49364
rect 29316 49308 31276 49364
rect 31332 49308 31342 49364
rect 13794 49196 13804 49252
rect 13860 49196 14812 49252
rect 14868 49196 19292 49252
rect 19348 49196 23212 49252
rect 23268 49196 23884 49252
rect 23940 49196 23950 49252
rect 27122 49196 27132 49252
rect 27188 49196 27916 49252
rect 27972 49196 27982 49252
rect 29922 49196 29932 49252
rect 29988 49196 42308 49252
rect 18386 49084 18396 49140
rect 18452 49084 19068 49140
rect 19124 49084 19134 49140
rect 20738 49084 20748 49140
rect 20804 49084 21756 49140
rect 21812 49084 21868 49140
rect 21924 49084 28812 49140
rect 28868 49084 28878 49140
rect 30370 49084 30380 49140
rect 30436 49084 31612 49140
rect 31668 49084 34524 49140
rect 34580 49084 34590 49140
rect 38994 49084 39004 49140
rect 39060 49084 39564 49140
rect 39620 49084 39630 49140
rect 42252 49028 42308 49196
rect 59200 49140 60000 49168
rect 43586 49084 43596 49140
rect 43652 49084 47740 49140
rect 47796 49084 47806 49140
rect 58258 49084 58268 49140
rect 58324 49084 60000 49140
rect 59200 49056 60000 49084
rect 13570 48972 13580 49028
rect 13636 48972 16604 49028
rect 16660 48972 16670 49028
rect 18946 48972 18956 49028
rect 19012 48972 20300 49028
rect 20356 48972 20366 49028
rect 21634 48972 21644 49028
rect 21700 48972 22876 49028
rect 22932 48972 22942 49028
rect 27010 48972 27020 49028
rect 27076 48972 27468 49028
rect 27524 48972 27534 49028
rect 28018 48972 28028 49028
rect 28084 48972 30044 49028
rect 30100 48972 30604 49028
rect 30660 48972 30670 49028
rect 33282 48972 33292 49028
rect 33348 48972 34076 49028
rect 34132 48972 34142 49028
rect 35522 48972 35532 49028
rect 35588 48972 37884 49028
rect 37940 48972 37950 49028
rect 38434 48972 38444 49028
rect 38500 48972 39452 49028
rect 39508 48972 39518 49028
rect 42242 48972 42252 49028
rect 42308 48972 42318 49028
rect 42802 48972 42812 49028
rect 42868 48972 43260 49028
rect 43316 48972 43326 49028
rect 19282 48860 19292 48916
rect 19348 48860 21532 48916
rect 21588 48860 21598 48916
rect 26852 48860 38668 48916
rect 42914 48860 42924 48916
rect 42980 48860 43932 48916
rect 43988 48860 43998 48916
rect 49074 48860 49084 48916
rect 49140 48860 50876 48916
rect 50932 48860 50942 48916
rect 26852 48804 26908 48860
rect 38612 48804 38668 48860
rect 16594 48748 16604 48804
rect 16660 48748 21308 48804
rect 21364 48748 21374 48804
rect 23174 48748 23212 48804
rect 23268 48748 23278 48804
rect 24322 48748 24332 48804
rect 24388 48748 26908 48804
rect 28578 48748 28588 48804
rect 28644 48748 30828 48804
rect 30884 48748 30894 48804
rect 31350 48748 31388 48804
rect 31444 48748 31454 48804
rect 33058 48748 33068 48804
rect 33124 48748 35644 48804
rect 35700 48748 36540 48804
rect 36596 48748 36606 48804
rect 38612 48748 39004 48804
rect 39060 48748 39070 48804
rect 42998 48748 43036 48804
rect 43092 48748 43102 48804
rect 43586 48748 43596 48804
rect 43652 48748 44156 48804
rect 44212 48748 44222 48804
rect 46050 48748 46060 48804
rect 46116 48748 47180 48804
rect 47236 48748 47516 48804
rect 47572 48748 47582 48804
rect 13906 48636 13916 48692
rect 13972 48636 16156 48692
rect 16212 48636 16222 48692
rect 22530 48636 22540 48692
rect 22596 48636 24556 48692
rect 24612 48636 24622 48692
rect 27318 48636 27356 48692
rect 27412 48636 27422 48692
rect 30258 48636 30268 48692
rect 30324 48636 30492 48692
rect 30548 48636 30558 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 22754 48524 22764 48580
rect 22820 48524 23324 48580
rect 23380 48524 23390 48580
rect 26114 48524 26124 48580
rect 26180 48524 30604 48580
rect 30660 48524 30670 48580
rect 40226 48524 40236 48580
rect 40292 48524 43932 48580
rect 43988 48524 43998 48580
rect 59200 48468 60000 48496
rect 21634 48412 21644 48468
rect 21700 48412 22876 48468
rect 22932 48412 22942 48468
rect 26450 48412 26460 48468
rect 26516 48412 26908 48468
rect 27122 48412 27132 48468
rect 27188 48412 27580 48468
rect 27636 48412 27646 48468
rect 32162 48412 32172 48468
rect 32228 48412 35420 48468
rect 35476 48412 35486 48468
rect 44930 48412 44940 48468
rect 44996 48412 49980 48468
rect 50036 48412 50988 48468
rect 51044 48412 51054 48468
rect 58146 48412 58156 48468
rect 58212 48412 60000 48468
rect 26852 48356 26908 48412
rect 59200 48384 60000 48412
rect 26852 48300 38556 48356
rect 38612 48300 38622 48356
rect 39778 48300 39788 48356
rect 39844 48300 42140 48356
rect 42196 48300 42206 48356
rect 42466 48300 42476 48356
rect 42532 48300 43148 48356
rect 43204 48300 44044 48356
rect 44100 48300 44604 48356
rect 44660 48300 44670 48356
rect 13346 48188 13356 48244
rect 13412 48188 14140 48244
rect 14196 48188 14206 48244
rect 22614 48188 22652 48244
rect 22708 48188 23548 48244
rect 23604 48188 23614 48244
rect 25890 48188 25900 48244
rect 25956 48188 26460 48244
rect 26516 48188 27580 48244
rect 27636 48188 27646 48244
rect 28018 48188 28028 48244
rect 28084 48188 28364 48244
rect 28420 48188 28924 48244
rect 28980 48188 28990 48244
rect 29922 48188 29932 48244
rect 29988 48188 30828 48244
rect 30884 48188 32060 48244
rect 32116 48188 32126 48244
rect 33842 48188 33852 48244
rect 33908 48188 34076 48244
rect 34132 48188 36540 48244
rect 36596 48188 36606 48244
rect 38322 48188 38332 48244
rect 38388 48188 39116 48244
rect 39172 48188 39182 48244
rect 39442 48188 39452 48244
rect 39508 48188 40012 48244
rect 40068 48188 40078 48244
rect 44930 48188 44940 48244
rect 44996 48188 45612 48244
rect 45668 48188 45678 48244
rect 15362 48076 15372 48132
rect 15428 48076 15708 48132
rect 15764 48076 16268 48132
rect 16324 48076 17164 48132
rect 17220 48076 17230 48132
rect 18470 48076 18508 48132
rect 18564 48076 18574 48132
rect 20738 48076 20748 48132
rect 20804 48076 25116 48132
rect 25172 48076 25182 48132
rect 25526 48076 25564 48132
rect 25620 48076 25630 48132
rect 20178 47964 20188 48020
rect 20244 47964 20748 48020
rect 20804 47964 20814 48020
rect 22306 47964 22316 48020
rect 22372 47964 23548 48020
rect 23604 47964 23614 48020
rect 24658 47964 24668 48020
rect 24724 47964 25676 48020
rect 25732 47964 25742 48020
rect 26852 47908 26908 48132
rect 26964 48076 26974 48132
rect 40226 48076 40236 48132
rect 40292 48076 41020 48132
rect 41076 48076 41086 48132
rect 40114 47964 40124 48020
rect 40180 47964 45388 48020
rect 45444 47964 45454 48020
rect 23986 47852 23996 47908
rect 24052 47852 26348 47908
rect 26404 47852 26908 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 17938 47740 17948 47796
rect 18004 47740 18844 47796
rect 18900 47740 18910 47796
rect 22866 47740 22876 47796
rect 22932 47740 33628 47796
rect 33684 47740 33694 47796
rect 22978 47628 22988 47684
rect 23044 47628 25676 47684
rect 25732 47628 25742 47684
rect 30146 47628 30156 47684
rect 30212 47628 33404 47684
rect 33460 47628 34300 47684
rect 34356 47628 36316 47684
rect 36372 47628 37436 47684
rect 37492 47628 37502 47684
rect 19618 47516 19628 47572
rect 19684 47516 21196 47572
rect 21252 47516 21262 47572
rect 22726 47516 22764 47572
rect 22820 47516 22830 47572
rect 27346 47516 27356 47572
rect 27412 47516 29932 47572
rect 29988 47516 29998 47572
rect 37650 47516 37660 47572
rect 37716 47516 40236 47572
rect 40292 47516 40302 47572
rect 49298 47516 49308 47572
rect 49364 47516 50652 47572
rect 50708 47516 50718 47572
rect 16706 47404 16716 47460
rect 16772 47404 19292 47460
rect 19348 47404 20636 47460
rect 20692 47404 20702 47460
rect 21522 47404 21532 47460
rect 21588 47404 22540 47460
rect 22596 47404 22606 47460
rect 24770 47404 24780 47460
rect 24836 47404 26124 47460
rect 26180 47404 26190 47460
rect 28130 47404 28140 47460
rect 28196 47404 29260 47460
rect 29316 47404 29326 47460
rect 29586 47404 29596 47460
rect 29652 47404 31164 47460
rect 31220 47404 31230 47460
rect 36530 47404 36540 47460
rect 36596 47404 37212 47460
rect 37268 47404 37278 47460
rect 46386 47404 46396 47460
rect 46452 47404 49532 47460
rect 49588 47404 50428 47460
rect 50484 47404 50494 47460
rect 53218 47404 53228 47460
rect 53284 47404 55580 47460
rect 55636 47404 55646 47460
rect 16716 47236 16772 47404
rect 17826 47292 17836 47348
rect 17892 47292 19740 47348
rect 19796 47292 19806 47348
rect 20514 47292 20524 47348
rect 20580 47292 25228 47348
rect 25284 47292 25294 47348
rect 27458 47292 27468 47348
rect 27524 47292 28252 47348
rect 28308 47292 28318 47348
rect 30818 47292 30828 47348
rect 30884 47292 31500 47348
rect 31556 47292 31566 47348
rect 38098 47292 38108 47348
rect 38164 47292 45500 47348
rect 45556 47292 45566 47348
rect 12450 47180 12460 47236
rect 12516 47180 15596 47236
rect 15652 47180 16772 47236
rect 17490 47180 17500 47236
rect 17556 47180 18396 47236
rect 18452 47180 18462 47236
rect 18610 47180 18620 47236
rect 18676 47180 18714 47236
rect 19394 47180 19404 47236
rect 19460 47180 20300 47236
rect 20356 47180 20366 47236
rect 20626 47180 20636 47236
rect 20692 47180 21196 47236
rect 21252 47180 21262 47236
rect 21634 47180 21644 47236
rect 21700 47180 22204 47236
rect 22260 47180 22270 47236
rect 22866 47180 22876 47236
rect 22932 47180 23324 47236
rect 23380 47180 23390 47236
rect 23482 47180 23492 47236
rect 23548 47180 24108 47236
rect 24164 47180 24174 47236
rect 27318 47180 27356 47236
rect 27412 47180 27422 47236
rect 31154 47180 31164 47236
rect 31220 47180 32620 47236
rect 32676 47180 32686 47236
rect 36306 47180 36316 47236
rect 36372 47180 37100 47236
rect 37156 47180 37166 47236
rect 38612 47180 39340 47236
rect 39396 47180 39406 47236
rect 18470 47068 18508 47124
rect 18564 47068 18574 47124
rect 19030 47068 19068 47124
rect 19124 47068 19134 47124
rect 19394 47068 19404 47124
rect 19460 47068 19628 47124
rect 19684 47068 19694 47124
rect 21298 47068 21308 47124
rect 21364 47068 23548 47124
rect 23604 47068 24220 47124
rect 24276 47068 24286 47124
rect 24994 47068 25004 47124
rect 25060 47068 26684 47124
rect 26740 47068 27468 47124
rect 27524 47068 28364 47124
rect 28420 47068 28430 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 38612 47012 38668 47180
rect 59200 47124 60000 47152
rect 39106 47068 39116 47124
rect 39172 47068 40012 47124
rect 40068 47068 40078 47124
rect 43474 47068 43484 47124
rect 43540 47068 45164 47124
rect 45220 47068 45230 47124
rect 57922 47068 57932 47124
rect 57988 47068 60000 47124
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 59200 47040 60000 47068
rect 13542 46956 13580 47012
rect 13636 46956 13646 47012
rect 16034 46956 16044 47012
rect 16100 46956 16604 47012
rect 16660 46956 17948 47012
rect 18004 46956 18014 47012
rect 18498 46956 18508 47012
rect 18564 46956 19292 47012
rect 19348 46956 19516 47012
rect 19572 46956 19582 47012
rect 23426 46956 23436 47012
rect 23492 46956 23548 47012
rect 23604 46956 23614 47012
rect 23772 46956 28028 47012
rect 28084 46956 28094 47012
rect 31266 46956 31276 47012
rect 31332 46956 38668 47012
rect 23772 46900 23828 46956
rect 16818 46844 16828 46900
rect 16884 46844 19628 46900
rect 19684 46844 20300 46900
rect 20356 46844 20366 46900
rect 22642 46844 22652 46900
rect 22708 46844 23324 46900
rect 23380 46844 23390 46900
rect 23762 46844 23772 46900
rect 23828 46844 23838 46900
rect 25330 46844 25340 46900
rect 25396 46844 25900 46900
rect 25956 46844 25966 46900
rect 39890 46844 39900 46900
rect 39956 46844 41020 46900
rect 41076 46844 41086 46900
rect 15026 46732 15036 46788
rect 15092 46732 18060 46788
rect 18116 46732 21308 46788
rect 21364 46732 21374 46788
rect 22978 46732 22988 46788
rect 23044 46732 23660 46788
rect 23716 46732 23726 46788
rect 23874 46732 23884 46788
rect 23940 46732 23978 46788
rect 24546 46732 24556 46788
rect 24612 46732 26796 46788
rect 26852 46732 26862 46788
rect 42018 46732 42028 46788
rect 42084 46732 44156 46788
rect 44212 46732 44222 46788
rect 46498 46732 46508 46788
rect 46564 46732 46732 46788
rect 46788 46732 46798 46788
rect 17826 46620 17836 46676
rect 17892 46620 18508 46676
rect 18564 46620 18574 46676
rect 19058 46620 19068 46676
rect 19124 46620 27020 46676
rect 27076 46620 27086 46676
rect 27234 46620 27244 46676
rect 27300 46620 28700 46676
rect 28756 46620 28766 46676
rect 30790 46620 30828 46676
rect 30884 46620 30894 46676
rect 41794 46620 41804 46676
rect 41860 46620 42588 46676
rect 42644 46620 42654 46676
rect 45378 46620 45388 46676
rect 45444 46620 46956 46676
rect 47012 46620 47022 46676
rect 49858 46620 49868 46676
rect 49924 46620 50652 46676
rect 50708 46620 50718 46676
rect 51314 46620 51324 46676
rect 51380 46620 53340 46676
rect 53396 46620 53406 46676
rect 8194 46508 8204 46564
rect 8260 46508 11228 46564
rect 11284 46508 11294 46564
rect 16258 46508 16268 46564
rect 16324 46508 17724 46564
rect 17780 46508 17790 46564
rect 21410 46508 21420 46564
rect 21476 46508 23212 46564
rect 23268 46508 24444 46564
rect 24500 46508 24510 46564
rect 27682 46508 27692 46564
rect 27748 46508 29036 46564
rect 29092 46508 29102 46564
rect 30482 46508 30492 46564
rect 30548 46508 31164 46564
rect 31220 46508 31230 46564
rect 48178 46508 48188 46564
rect 48244 46508 49532 46564
rect 49588 46508 49598 46564
rect 51650 46508 51660 46564
rect 51716 46508 53116 46564
rect 53172 46508 53182 46564
rect 9874 46396 9884 46452
rect 9940 46396 12460 46452
rect 12516 46396 12684 46452
rect 12740 46396 12750 46452
rect 13010 46396 13020 46452
rect 13076 46396 14140 46452
rect 14196 46396 14206 46452
rect 16482 46396 16492 46452
rect 16548 46396 17388 46452
rect 17444 46396 17454 46452
rect 20402 46396 20412 46452
rect 20468 46396 20748 46452
rect 20804 46396 20814 46452
rect 22082 46396 22092 46452
rect 22148 46396 22158 46452
rect 22530 46396 22540 46452
rect 22596 46396 25788 46452
rect 25844 46396 26460 46452
rect 26516 46396 26526 46452
rect 26758 46396 26796 46452
rect 26852 46396 26862 46452
rect 22092 46340 22148 46396
rect 22092 46284 22428 46340
rect 22484 46284 22494 46340
rect 26562 46284 26572 46340
rect 26628 46284 27916 46340
rect 27972 46284 27982 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 16706 46172 16716 46228
rect 16772 46172 18284 46228
rect 18340 46172 18732 46228
rect 18788 46172 18798 46228
rect 19954 46172 19964 46228
rect 20020 46172 20860 46228
rect 20916 46172 20926 46228
rect 21970 46172 21980 46228
rect 22036 46172 23884 46228
rect 23940 46172 23950 46228
rect 27766 46172 27804 46228
rect 27860 46172 27870 46228
rect 27990 46172 28028 46228
rect 28084 46172 28094 46228
rect 12338 46060 12348 46116
rect 12404 46060 13692 46116
rect 13748 46060 14588 46116
rect 14644 46060 14654 46116
rect 17938 46060 17948 46116
rect 18004 46060 18014 46116
rect 18498 46060 18508 46116
rect 18564 46060 18844 46116
rect 18900 46060 20636 46116
rect 20692 46060 20702 46116
rect 23090 46060 23100 46116
rect 23156 46060 23436 46116
rect 23492 46060 23502 46116
rect 26674 46060 26684 46116
rect 26740 46060 29708 46116
rect 29764 46060 29774 46116
rect 29922 46060 29932 46116
rect 29988 46060 31500 46116
rect 31556 46060 31566 46116
rect 35858 46060 35868 46116
rect 35924 46060 45052 46116
rect 45108 46060 45118 46116
rect 17948 46004 18004 46060
rect 12450 45948 12460 46004
rect 12516 45948 14028 46004
rect 14084 45948 14094 46004
rect 14354 45948 14364 46004
rect 14420 45948 16828 46004
rect 16884 45948 16894 46004
rect 17490 45948 17500 46004
rect 17556 45948 18004 46004
rect 18274 45948 18284 46004
rect 18340 45948 27692 46004
rect 27748 45948 27758 46004
rect 32498 45948 32508 46004
rect 32564 45948 34300 46004
rect 34356 45948 34366 46004
rect 34626 45948 34636 46004
rect 34692 45948 35196 46004
rect 35252 45948 35262 46004
rect 14242 45836 14252 45892
rect 14308 45836 14924 45892
rect 14980 45836 14990 45892
rect 15586 45836 15596 45892
rect 15652 45836 15932 45892
rect 15988 45836 16268 45892
rect 16324 45836 16334 45892
rect 16930 45836 16940 45892
rect 16996 45836 17724 45892
rect 17780 45836 17790 45892
rect 17938 45836 17948 45892
rect 18004 45836 18620 45892
rect 18676 45836 18686 45892
rect 18834 45836 18844 45892
rect 18900 45836 20076 45892
rect 20132 45836 21868 45892
rect 21924 45836 21934 45892
rect 25666 45836 25676 45892
rect 25732 45836 27020 45892
rect 27076 45836 27524 45892
rect 28354 45836 28364 45892
rect 28420 45836 30156 45892
rect 30212 45836 31612 45892
rect 31668 45836 31678 45892
rect 32834 45836 32844 45892
rect 32900 45836 33516 45892
rect 33572 45836 35084 45892
rect 35140 45836 35150 45892
rect 43810 45836 43820 45892
rect 43876 45836 46844 45892
rect 46900 45836 46910 45892
rect 50306 45836 50316 45892
rect 50372 45836 51660 45892
rect 51716 45836 52444 45892
rect 52500 45836 52510 45892
rect 27468 45780 27524 45836
rect 16034 45724 16044 45780
rect 16100 45724 25228 45780
rect 25284 45724 25294 45780
rect 27468 45724 29260 45780
rect 29316 45724 29326 45780
rect 30034 45724 30044 45780
rect 30100 45724 31164 45780
rect 31220 45724 31230 45780
rect 31826 45724 31836 45780
rect 31892 45724 33740 45780
rect 33796 45724 34524 45780
rect 34580 45724 34590 45780
rect 39442 45724 39452 45780
rect 39508 45724 43708 45780
rect 43764 45724 43774 45780
rect 13458 45612 13468 45668
rect 13524 45612 14252 45668
rect 14308 45612 14812 45668
rect 14868 45612 14878 45668
rect 15586 45612 15596 45668
rect 15652 45612 18844 45668
rect 18900 45612 18910 45668
rect 19058 45612 19068 45668
rect 19124 45612 19516 45668
rect 19572 45612 20300 45668
rect 20356 45612 23548 45668
rect 28018 45612 28028 45668
rect 28084 45612 28140 45668
rect 28196 45612 28206 45668
rect 29698 45612 29708 45668
rect 29764 45612 30604 45668
rect 30660 45612 30670 45668
rect 23492 45556 23548 45612
rect 12786 45500 12796 45556
rect 12852 45500 16492 45556
rect 16548 45500 16558 45556
rect 23492 45500 24444 45556
rect 24500 45500 26908 45556
rect 26964 45500 26974 45556
rect 44146 45500 44156 45556
rect 44212 45500 44940 45556
rect 44996 45500 45006 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 15474 45388 15484 45444
rect 15540 45388 17388 45444
rect 17444 45388 17454 45444
rect 25778 45388 25788 45444
rect 25844 45388 26572 45444
rect 26628 45388 26638 45444
rect 31826 45388 31836 45444
rect 31892 45388 32844 45444
rect 32900 45388 32910 45444
rect 10546 45276 10556 45332
rect 10612 45276 14364 45332
rect 14420 45276 14924 45332
rect 14980 45276 14990 45332
rect 15092 45276 18284 45332
rect 18340 45276 18350 45332
rect 18732 45276 18844 45332
rect 18900 45276 19516 45332
rect 19572 45276 19582 45332
rect 22194 45276 22204 45332
rect 22260 45276 25340 45332
rect 25396 45276 25406 45332
rect 26114 45276 26124 45332
rect 26180 45276 26684 45332
rect 26740 45276 26750 45332
rect 41234 45276 41244 45332
rect 41300 45276 42700 45332
rect 42756 45276 42766 45332
rect 15092 45220 15148 45276
rect 18732 45220 18788 45276
rect 8082 45164 8092 45220
rect 8148 45164 15148 45220
rect 15362 45164 15372 45220
rect 15428 45164 16716 45220
rect 16772 45164 16782 45220
rect 17042 45164 17052 45220
rect 17108 45164 18788 45220
rect 19058 45164 19068 45220
rect 19124 45164 24444 45220
rect 24500 45164 27132 45220
rect 27188 45164 27198 45220
rect 37986 45164 37996 45220
rect 38052 45164 40908 45220
rect 40964 45164 40974 45220
rect 11116 45052 15148 45108
rect 17714 45052 17724 45108
rect 17780 45052 19852 45108
rect 19908 45052 19918 45108
rect 22530 45052 22540 45108
rect 22596 45052 24332 45108
rect 24388 45052 26236 45108
rect 26292 45052 26302 45108
rect 26852 45052 27468 45108
rect 27524 45052 27534 45108
rect 28550 45052 28588 45108
rect 28644 45052 28654 45108
rect 34374 45052 34412 45108
rect 34468 45052 34478 45108
rect 37874 45052 37884 45108
rect 37940 45052 38668 45108
rect 39442 45052 39452 45108
rect 39508 45052 42252 45108
rect 42308 45052 42318 45108
rect 11116 44996 11172 45052
rect 15092 44996 15148 45052
rect 11106 44940 11116 44996
rect 11172 44940 11182 44996
rect 14466 44940 14476 44996
rect 14532 44940 14542 44996
rect 15092 44940 16044 44996
rect 16100 44940 16110 44996
rect 16258 44940 16268 44996
rect 16324 44940 18172 44996
rect 18228 44940 18238 44996
rect 18396 44940 22092 44996
rect 22148 44940 22652 44996
rect 22708 44940 22718 44996
rect 26786 44940 26796 44996
rect 26852 44940 26908 45052
rect 38612 44996 38668 45052
rect 27468 44940 28028 44996
rect 28084 44940 28094 44996
rect 30930 44940 30940 44996
rect 30996 44940 31948 44996
rect 32004 44940 32014 44996
rect 34178 44940 34188 44996
rect 34244 44940 35196 44996
rect 35252 44940 35262 44996
rect 38612 44940 38948 44996
rect 39778 44940 39788 44996
rect 39844 44940 41244 44996
rect 41300 44940 41310 44996
rect 42354 44940 42364 44996
rect 42420 44940 47404 44996
rect 47460 44940 47470 44996
rect 14476 44772 14532 44940
rect 18396 44884 18452 44940
rect 27468 44884 27524 44940
rect 38892 44884 38948 44940
rect 16930 44828 16940 44884
rect 16996 44828 18452 44884
rect 19954 44828 19964 44884
rect 20020 44828 23436 44884
rect 23492 44772 23548 44884
rect 23650 44828 23660 44884
rect 23716 44828 25004 44884
rect 25060 44828 25070 44884
rect 25442 44828 25452 44884
rect 25508 44828 25676 44884
rect 25732 44828 27524 44884
rect 28130 44828 28140 44884
rect 28196 44828 31388 44884
rect 31444 44828 31454 44884
rect 34972 44828 38668 44884
rect 38892 44828 39116 44884
rect 39172 44828 39182 44884
rect 50082 44828 50092 44884
rect 50148 44828 50876 44884
rect 50932 44828 50942 44884
rect 34972 44772 35028 44828
rect 14476 44716 23100 44772
rect 23156 44716 23166 44772
rect 23492 44716 28588 44772
rect 28644 44716 28654 44772
rect 29698 44716 29708 44772
rect 29764 44716 35028 44772
rect 38612 44772 38668 44828
rect 38612 44716 38780 44772
rect 38836 44716 38846 44772
rect 47730 44716 47740 44772
rect 47796 44716 49532 44772
rect 49588 44716 49598 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 13010 44604 13020 44660
rect 13076 44604 13692 44660
rect 13748 44604 17052 44660
rect 17108 44604 17118 44660
rect 17602 44604 17612 44660
rect 17668 44604 22764 44660
rect 22820 44604 22830 44660
rect 26898 44604 26908 44660
rect 26964 44604 34300 44660
rect 34356 44604 34366 44660
rect 14130 44492 14140 44548
rect 14196 44492 15036 44548
rect 15092 44492 15102 44548
rect 15782 44492 15820 44548
rect 15876 44492 15886 44548
rect 17042 44492 17052 44548
rect 17108 44492 17388 44548
rect 17444 44492 17454 44548
rect 19282 44492 19292 44548
rect 19348 44492 20524 44548
rect 20580 44492 20590 44548
rect 21858 44492 21868 44548
rect 21924 44492 23660 44548
rect 23716 44492 23726 44548
rect 26852 44492 30492 44548
rect 30548 44492 30558 44548
rect 37314 44492 37324 44548
rect 37380 44492 46172 44548
rect 46228 44492 46238 44548
rect 26852 44436 26908 44492
rect 14354 44380 14364 44436
rect 14420 44380 14588 44436
rect 14644 44380 15372 44436
rect 15428 44380 15438 44436
rect 15708 44380 16268 44436
rect 16324 44380 16334 44436
rect 16706 44380 16716 44436
rect 16772 44380 26908 44436
rect 28578 44380 28588 44436
rect 28644 44380 29484 44436
rect 29540 44380 29550 44436
rect 38658 44380 38668 44436
rect 38724 44380 39676 44436
rect 39732 44380 40460 44436
rect 40516 44380 40526 44436
rect 15708 44324 15764 44380
rect 10098 44268 10108 44324
rect 10164 44268 10892 44324
rect 10948 44268 10958 44324
rect 12002 44268 12012 44324
rect 12068 44268 13580 44324
rect 13636 44268 15764 44324
rect 15922 44268 15932 44324
rect 15988 44268 17052 44324
rect 17108 44268 17836 44324
rect 17892 44268 17902 44324
rect 19058 44268 19068 44324
rect 19124 44268 19516 44324
rect 19572 44268 21308 44324
rect 21364 44268 21374 44324
rect 21746 44268 21756 44324
rect 21812 44268 22428 44324
rect 22484 44268 22494 44324
rect 23650 44268 23660 44324
rect 23716 44268 23726 44324
rect 24434 44268 24444 44324
rect 24500 44268 25340 44324
rect 25396 44268 25406 44324
rect 26002 44268 26012 44324
rect 26068 44268 28252 44324
rect 28308 44268 29932 44324
rect 29988 44268 29998 44324
rect 30594 44268 30604 44324
rect 30660 44268 30940 44324
rect 30996 44268 32284 44324
rect 32340 44268 32350 44324
rect 35298 44268 35308 44324
rect 35364 44268 36988 44324
rect 37044 44268 37054 44324
rect 38770 44268 38780 44324
rect 38836 44268 45948 44324
rect 46004 44268 46396 44324
rect 46452 44268 46462 44324
rect 46834 44268 46844 44324
rect 46900 44268 47516 44324
rect 47572 44268 47582 44324
rect 52994 44268 53004 44324
rect 53060 44268 55580 44324
rect 55636 44268 55646 44324
rect 23660 44212 23716 44268
rect 17490 44156 17500 44212
rect 17556 44156 22652 44212
rect 22708 44156 23324 44212
rect 23380 44156 23390 44212
rect 23660 44156 29708 44212
rect 29764 44156 29774 44212
rect 38612 44156 39228 44212
rect 39284 44156 40124 44212
rect 40180 44156 40628 44212
rect 41346 44156 41356 44212
rect 41412 44156 41916 44212
rect 41972 44156 42700 44212
rect 42756 44156 42766 44212
rect 10322 44044 10332 44100
rect 10388 44044 11788 44100
rect 16482 44044 16492 44100
rect 16548 44044 17724 44100
rect 17780 44044 17790 44100
rect 17938 44044 17948 44100
rect 18004 44044 18060 44100
rect 18116 44044 19628 44100
rect 19684 44044 19694 44100
rect 22082 44044 22092 44100
rect 22148 44044 23548 44100
rect 23604 44044 23614 44100
rect 11732 43988 11788 44044
rect 11732 43932 12572 43988
rect 12628 43932 18844 43988
rect 18900 43932 18910 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 38612 43876 38668 44156
rect 40572 44100 40628 44156
rect 40572 44044 41020 44100
rect 41076 44044 41086 44100
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 10434 43820 10444 43876
rect 10500 43820 11228 43876
rect 11284 43820 11294 43876
rect 19282 43820 19292 43876
rect 19348 43820 19358 43876
rect 21746 43820 21756 43876
rect 21812 43820 38332 43876
rect 38388 43820 38668 43876
rect 15708 43708 16268 43764
rect 16324 43708 16334 43764
rect 18694 43708 18732 43764
rect 18788 43708 18798 43764
rect 15708 43540 15764 43708
rect 16146 43596 16156 43652
rect 16212 43596 16380 43652
rect 16436 43596 16446 43652
rect 16594 43596 16604 43652
rect 16660 43596 17612 43652
rect 17668 43596 17678 43652
rect 16380 43540 16436 43596
rect 19292 43540 19348 43820
rect 59200 43764 60000 43792
rect 57922 43708 57932 43764
rect 57988 43708 60000 43764
rect 59200 43680 60000 43708
rect 20962 43596 20972 43652
rect 21028 43596 23884 43652
rect 23940 43596 23950 43652
rect 26898 43596 26908 43652
rect 26964 43596 38668 43652
rect 48290 43596 48300 43652
rect 48356 43596 49756 43652
rect 49812 43596 49822 43652
rect 9986 43484 9996 43540
rect 10052 43484 10444 43540
rect 10500 43484 10780 43540
rect 10836 43484 12460 43540
rect 12516 43484 12526 43540
rect 15670 43484 15708 43540
rect 15764 43484 15774 43540
rect 16380 43484 16940 43540
rect 16996 43484 17724 43540
rect 17780 43484 17790 43540
rect 18722 43484 18732 43540
rect 18788 43484 19348 43540
rect 23314 43484 23324 43540
rect 23380 43484 25228 43540
rect 25284 43484 25294 43540
rect 26310 43484 26348 43540
rect 26404 43484 26414 43540
rect 27570 43484 27580 43540
rect 27636 43484 32284 43540
rect 32340 43484 32350 43540
rect 33842 43484 33852 43540
rect 33908 43484 34748 43540
rect 34804 43484 34814 43540
rect 36306 43484 36316 43540
rect 36372 43484 38108 43540
rect 38164 43484 38174 43540
rect 34748 43428 34804 43484
rect 10892 43372 19292 43428
rect 19348 43372 19628 43428
rect 19684 43372 19694 43428
rect 22978 43372 22988 43428
rect 23044 43372 25564 43428
rect 25620 43372 25630 43428
rect 30482 43372 30492 43428
rect 30548 43372 31948 43428
rect 32004 43372 32620 43428
rect 32676 43372 32686 43428
rect 34748 43372 37548 43428
rect 37604 43372 37884 43428
rect 37940 43372 37950 43428
rect 10892 43316 10948 43372
rect 38612 43316 38668 43596
rect 51090 43484 51100 43540
rect 51156 43484 52332 43540
rect 52388 43484 52398 43540
rect 50642 43372 50652 43428
rect 50708 43372 52444 43428
rect 52500 43372 52510 43428
rect 10882 43260 10892 43316
rect 10948 43260 10958 43316
rect 11554 43260 11564 43316
rect 11620 43260 13020 43316
rect 13076 43260 13086 43316
rect 13682 43260 13692 43316
rect 13748 43260 15484 43316
rect 15540 43260 15550 43316
rect 16370 43260 16380 43316
rect 16436 43260 18396 43316
rect 18452 43260 18732 43316
rect 18788 43260 18798 43316
rect 19842 43260 19852 43316
rect 19908 43260 25452 43316
rect 25508 43260 25518 43316
rect 26674 43260 26684 43316
rect 26740 43260 27580 43316
rect 27636 43260 27646 43316
rect 28102 43260 28140 43316
rect 28196 43260 28206 43316
rect 38612 43260 39228 43316
rect 39284 43260 39294 43316
rect 43138 43260 43148 43316
rect 43204 43260 45276 43316
rect 45332 43260 45342 43316
rect 49858 43260 49868 43316
rect 49924 43260 50876 43316
rect 50932 43260 51212 43316
rect 51268 43260 51278 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 15922 43036 15932 43092
rect 15988 43036 26572 43092
rect 26628 43036 27580 43092
rect 27636 43036 28476 43092
rect 28532 43036 28542 43092
rect 34262 43036 34300 43092
rect 34356 43036 34972 43092
rect 35028 43036 35038 43092
rect 38668 42980 38724 43260
rect 21298 42924 21308 42980
rect 21364 42924 22876 42980
rect 22932 42924 23268 42980
rect 23426 42924 23436 42980
rect 23492 42924 26908 42980
rect 27010 42924 27020 42980
rect 27076 42924 28196 42980
rect 37314 42924 37324 42980
rect 37380 42924 37884 42980
rect 37940 42924 37950 42980
rect 38658 42924 38668 42980
rect 38724 42924 38734 42980
rect 23212 42868 23268 42924
rect 26852 42868 26908 42924
rect 28140 42868 28196 42924
rect 16818 42812 16828 42868
rect 16884 42812 17388 42868
rect 17444 42812 17454 42868
rect 18162 42812 18172 42868
rect 18228 42812 21644 42868
rect 21700 42812 21710 42868
rect 23212 42812 24724 42868
rect 26852 42812 27468 42868
rect 27524 42812 27534 42868
rect 28130 42812 28140 42868
rect 28196 42812 30604 42868
rect 30660 42812 30670 42868
rect 34290 42812 34300 42868
rect 34356 42812 34860 42868
rect 34916 42812 35868 42868
rect 35924 42812 35934 42868
rect 43138 42812 43148 42868
rect 43204 42812 44940 42868
rect 44996 42812 45006 42868
rect 17388 42756 17444 42812
rect 24668 42756 24724 42812
rect 17388 42700 18284 42756
rect 18340 42700 18350 42756
rect 18806 42700 18844 42756
rect 18900 42700 18910 42756
rect 19058 42700 19068 42756
rect 19124 42700 19628 42756
rect 19684 42700 19694 42756
rect 19852 42700 21756 42756
rect 21812 42700 24220 42756
rect 24276 42700 24286 42756
rect 24658 42700 24668 42756
rect 24724 42700 24734 42756
rect 24882 42700 24892 42756
rect 24948 42700 30716 42756
rect 30772 42700 30782 42756
rect 38546 42700 38556 42756
rect 38612 42700 39004 42756
rect 39060 42700 39070 42756
rect 39890 42700 39900 42756
rect 39956 42700 42028 42756
rect 42084 42700 42094 42756
rect 50082 42700 50092 42756
rect 50148 42700 50764 42756
rect 50820 42700 50830 42756
rect 51762 42700 51772 42756
rect 51828 42700 55580 42756
rect 55636 42700 55646 42756
rect 19852 42644 19908 42700
rect 15586 42588 15596 42644
rect 15652 42588 16604 42644
rect 16660 42588 16670 42644
rect 17378 42588 17388 42644
rect 17444 42588 19908 42644
rect 20290 42588 20300 42644
rect 20356 42588 23660 42644
rect 23716 42588 23726 42644
rect 25666 42588 25676 42644
rect 25732 42588 27020 42644
rect 27076 42588 27086 42644
rect 28102 42588 28140 42644
rect 28196 42588 28206 42644
rect 30370 42588 30380 42644
rect 30436 42588 31388 42644
rect 31444 42588 31454 42644
rect 35634 42588 35644 42644
rect 35700 42588 38668 42644
rect 38612 42532 38668 42588
rect 12450 42476 12460 42532
rect 12516 42476 13580 42532
rect 13636 42476 13646 42532
rect 19730 42476 19740 42532
rect 19796 42476 20636 42532
rect 20692 42476 20702 42532
rect 20850 42476 20860 42532
rect 20916 42476 26124 42532
rect 26180 42476 26190 42532
rect 27458 42476 27468 42532
rect 27524 42476 28588 42532
rect 28644 42476 28654 42532
rect 31574 42476 31612 42532
rect 31668 42476 31678 42532
rect 38612 42476 43820 42532
rect 43876 42476 44828 42532
rect 44884 42476 44894 42532
rect 45042 42476 45052 42532
rect 45108 42476 45276 42532
rect 45332 42476 45612 42532
rect 45668 42476 45678 42532
rect 23538 42364 23548 42420
rect 23604 42364 25228 42420
rect 25284 42364 25294 42420
rect 26002 42364 26012 42420
rect 26068 42364 27020 42420
rect 27076 42364 27132 42420
rect 27188 42364 27198 42420
rect 27794 42364 27804 42420
rect 27860 42364 32172 42420
rect 32228 42364 32238 42420
rect 35298 42364 35308 42420
rect 35364 42364 35756 42420
rect 35812 42364 35822 42420
rect 41234 42364 41244 42420
rect 41300 42364 42140 42420
rect 42196 42364 43260 42420
rect 43316 42364 43326 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 18274 42252 18284 42308
rect 18340 42252 18732 42308
rect 18788 42252 18798 42308
rect 18946 42252 18956 42308
rect 19012 42252 19628 42308
rect 19684 42252 19694 42308
rect 20514 42252 20524 42308
rect 20580 42252 20590 42308
rect 20962 42252 20972 42308
rect 21028 42252 24556 42308
rect 24612 42252 24622 42308
rect 25554 42252 25564 42308
rect 25620 42252 26796 42308
rect 26852 42252 26862 42308
rect 27458 42252 27468 42308
rect 27524 42252 27580 42308
rect 27636 42252 27646 42308
rect 34262 42252 34300 42308
rect 34356 42252 34366 42308
rect 20524 42196 20580 42252
rect 15250 42140 15260 42196
rect 15316 42140 15354 42196
rect 16146 42140 16156 42196
rect 16212 42140 20580 42196
rect 21410 42140 21420 42196
rect 21476 42140 21644 42196
rect 21700 42140 22876 42196
rect 22932 42140 22942 42196
rect 23538 42140 23548 42196
rect 23604 42140 27356 42196
rect 27412 42140 27422 42196
rect 34738 42140 34748 42196
rect 34804 42140 35980 42196
rect 36036 42140 36046 42196
rect 38658 42140 38668 42196
rect 38724 42140 39676 42196
rect 39732 42140 40236 42196
rect 40292 42140 40302 42196
rect 47170 42140 47180 42196
rect 47236 42140 49196 42196
rect 49252 42140 49262 42196
rect 13234 42028 13244 42084
rect 13300 42028 14252 42084
rect 14308 42028 14588 42084
rect 14644 42028 14654 42084
rect 15026 42028 15036 42084
rect 15092 42028 19852 42084
rect 19908 42028 19918 42084
rect 20076 42028 22988 42084
rect 23044 42028 23054 42084
rect 23650 42028 23660 42084
rect 23716 42028 25452 42084
rect 25508 42028 25518 42084
rect 26534 42028 26572 42084
rect 26628 42028 26638 42084
rect 26786 42028 26796 42084
rect 26852 42028 30940 42084
rect 30996 42028 31006 42084
rect 33730 42028 33740 42084
rect 33796 42028 34412 42084
rect 34468 42028 34478 42084
rect 20076 41972 20132 42028
rect 13906 41916 13916 41972
rect 13972 41916 15260 41972
rect 15316 41916 15708 41972
rect 15764 41916 15774 41972
rect 16034 41916 16044 41972
rect 16100 41916 17388 41972
rect 17444 41916 17454 41972
rect 18386 41916 18396 41972
rect 18452 41916 20132 41972
rect 22642 41916 22652 41972
rect 22708 41916 24612 41972
rect 24770 41916 24780 41972
rect 24836 41916 26012 41972
rect 26068 41916 26078 41972
rect 27906 41916 27916 41972
rect 27972 41916 30268 41972
rect 30324 41916 30334 41972
rect 34626 41916 34636 41972
rect 34692 41916 35308 41972
rect 35364 41916 35374 41972
rect 46834 41916 46844 41972
rect 46900 41916 48412 41972
rect 48468 41916 48478 41972
rect 24556 41860 24612 41916
rect 19170 41804 19180 41860
rect 19236 41804 23212 41860
rect 23268 41804 23278 41860
rect 24556 41804 26348 41860
rect 26404 41804 26414 41860
rect 26674 41804 26684 41860
rect 26740 41804 27860 41860
rect 28662 41804 28700 41860
rect 28756 41804 28766 41860
rect 32498 41804 32508 41860
rect 32564 41804 33180 41860
rect 33236 41804 34300 41860
rect 34356 41804 34366 41860
rect 8866 41692 8876 41748
rect 8932 41692 14476 41748
rect 14532 41692 15260 41748
rect 15316 41692 15326 41748
rect 20402 41692 20412 41748
rect 20468 41692 23772 41748
rect 23828 41692 23838 41748
rect 24546 41692 24556 41748
rect 24612 41692 24622 41748
rect 15138 41580 15148 41636
rect 15204 41580 15260 41636
rect 15316 41580 15326 41636
rect 16034 41580 16044 41636
rect 16100 41580 20972 41636
rect 21028 41580 21038 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 24556 41524 24612 41692
rect 27804 41636 27860 41804
rect 59200 41748 60000 41776
rect 28018 41692 28028 41748
rect 28084 41692 29260 41748
rect 29316 41692 29326 41748
rect 39890 41692 39900 41748
rect 39956 41692 41020 41748
rect 41076 41692 42476 41748
rect 42532 41692 42542 41748
rect 44482 41692 44492 41748
rect 44548 41692 45836 41748
rect 45892 41692 47404 41748
rect 47460 41692 47470 41748
rect 57922 41692 57932 41748
rect 57988 41692 60000 41748
rect 59200 41664 60000 41692
rect 27804 41580 33516 41636
rect 33572 41580 33582 41636
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 11778 41468 11788 41524
rect 11844 41468 12684 41524
rect 12740 41468 12750 41524
rect 16146 41468 16156 41524
rect 16212 41468 18340 41524
rect 24556 41468 29148 41524
rect 29204 41468 29214 41524
rect 18284 41412 18340 41468
rect 14802 41356 14812 41412
rect 14868 41356 17276 41412
rect 17332 41356 17342 41412
rect 18274 41356 18284 41412
rect 18340 41356 18844 41412
rect 18900 41356 18910 41412
rect 19394 41356 19404 41412
rect 19460 41356 19964 41412
rect 20020 41356 21532 41412
rect 21588 41356 21598 41412
rect 23986 41356 23996 41412
rect 24052 41356 25228 41412
rect 25284 41356 25294 41412
rect 26534 41356 26572 41412
rect 26628 41356 26638 41412
rect 28130 41356 28140 41412
rect 28196 41356 32172 41412
rect 32228 41356 32238 41412
rect 1698 41244 1708 41300
rect 1764 41244 1774 41300
rect 10210 41244 10220 41300
rect 10276 41244 11004 41300
rect 11060 41244 11070 41300
rect 14578 41244 14588 41300
rect 14644 41244 15260 41300
rect 15316 41244 21980 41300
rect 22036 41244 22046 41300
rect 26982 41244 27020 41300
rect 27076 41244 27086 41300
rect 27570 41244 27580 41300
rect 27636 41244 28700 41300
rect 28756 41244 28766 41300
rect 32386 41244 32396 41300
rect 32452 41244 33516 41300
rect 33572 41244 33582 41300
rect 45154 41244 45164 41300
rect 45220 41244 45948 41300
rect 46004 41244 46014 41300
rect 0 41076 800 41104
rect 1708 41076 1764 41244
rect 9650 41132 9660 41188
rect 9716 41132 12348 41188
rect 12404 41132 12414 41188
rect 17266 41132 17276 41188
rect 17332 41132 25228 41188
rect 25284 41132 25294 41188
rect 27794 41132 27804 41188
rect 27860 41132 28028 41188
rect 28084 41132 28094 41188
rect 50418 41132 50428 41188
rect 50484 41132 55580 41188
rect 55636 41132 55646 41188
rect 0 41020 1764 41076
rect 12674 41020 12684 41076
rect 12740 41020 18396 41076
rect 18452 41020 19740 41076
rect 19796 41020 19806 41076
rect 21522 41020 21532 41076
rect 21588 41020 22428 41076
rect 22484 41020 22494 41076
rect 34402 41020 34412 41076
rect 34468 41020 35084 41076
rect 35140 41020 35150 41076
rect 0 40992 800 41020
rect 8754 40908 8764 40964
rect 8820 40908 9772 40964
rect 9828 40908 9838 40964
rect 12002 40908 12012 40964
rect 12068 40908 18060 40964
rect 18116 40908 18620 40964
rect 18676 40908 19516 40964
rect 19572 40908 19582 40964
rect 20290 40908 20300 40964
rect 20356 40908 21196 40964
rect 21252 40908 21262 40964
rect 31602 40908 31612 40964
rect 31668 40908 39564 40964
rect 39620 40908 39630 40964
rect 48066 40908 48076 40964
rect 48132 40908 49532 40964
rect 49588 40908 49598 40964
rect 22754 40796 22764 40852
rect 22820 40796 26124 40852
rect 26180 40796 26190 40852
rect 29138 40796 29148 40852
rect 29204 40796 30940 40852
rect 30996 40796 31006 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 12002 40684 12012 40740
rect 12068 40684 13468 40740
rect 13524 40684 15708 40740
rect 15764 40684 16716 40740
rect 16772 40684 16782 40740
rect 20710 40684 20748 40740
rect 20804 40684 20814 40740
rect 26226 40684 26236 40740
rect 26292 40684 33292 40740
rect 33348 40684 33358 40740
rect 10658 40572 10668 40628
rect 10724 40572 13356 40628
rect 13412 40572 13422 40628
rect 18946 40572 18956 40628
rect 19012 40572 22316 40628
rect 22372 40572 22988 40628
rect 23044 40572 23054 40628
rect 29362 40572 29372 40628
rect 29428 40572 29820 40628
rect 29876 40572 29886 40628
rect 31490 40572 31500 40628
rect 31556 40572 32172 40628
rect 32228 40572 33180 40628
rect 33236 40572 33246 40628
rect 13234 40460 13244 40516
rect 13300 40460 15148 40516
rect 15204 40460 16268 40516
rect 16324 40460 16334 40516
rect 16482 40460 16492 40516
rect 16548 40460 17724 40516
rect 17780 40460 17790 40516
rect 17938 40460 17948 40516
rect 18004 40460 18732 40516
rect 18788 40460 18798 40516
rect 19516 40460 24108 40516
rect 24164 40460 24174 40516
rect 24546 40460 24556 40516
rect 24612 40460 25340 40516
rect 25396 40460 25406 40516
rect 26786 40460 26796 40516
rect 26852 40460 28476 40516
rect 28532 40460 28542 40516
rect 33506 40460 33516 40516
rect 33572 40460 34300 40516
rect 34356 40460 34366 40516
rect 39442 40460 39452 40516
rect 39508 40460 39788 40516
rect 39844 40460 41356 40516
rect 41412 40460 42028 40516
rect 42084 40460 42094 40516
rect 16268 40404 16324 40460
rect 19516 40404 19572 40460
rect 59200 40404 60000 40432
rect 9762 40348 9772 40404
rect 9828 40348 11004 40404
rect 11060 40348 11070 40404
rect 11330 40348 11340 40404
rect 11396 40348 15036 40404
rect 15092 40348 15484 40404
rect 15540 40348 15550 40404
rect 16268 40348 17500 40404
rect 17556 40348 17566 40404
rect 19506 40348 19516 40404
rect 19572 40348 19582 40404
rect 19842 40348 19852 40404
rect 19908 40348 20524 40404
rect 20580 40348 20590 40404
rect 22418 40348 22428 40404
rect 22484 40348 27916 40404
rect 27972 40348 27982 40404
rect 29596 40348 34076 40404
rect 34132 40348 34142 40404
rect 39554 40348 39564 40404
rect 39620 40348 41580 40404
rect 41636 40348 41646 40404
rect 47842 40348 47852 40404
rect 47908 40348 49084 40404
rect 49140 40348 49150 40404
rect 57922 40348 57932 40404
rect 57988 40348 60000 40404
rect 11004 40292 11060 40348
rect 11004 40236 12684 40292
rect 12740 40236 12750 40292
rect 13458 40236 13468 40292
rect 13524 40236 14812 40292
rect 14868 40236 14878 40292
rect 15586 40236 15596 40292
rect 15652 40236 20356 40292
rect 20626 40236 20636 40292
rect 20692 40236 21532 40292
rect 21588 40236 21598 40292
rect 12684 40180 12740 40236
rect 20300 40180 20356 40236
rect 29596 40180 29652 40348
rect 59200 40320 60000 40348
rect 34850 40236 34860 40292
rect 34916 40236 36316 40292
rect 36372 40236 36382 40292
rect 43810 40236 43820 40292
rect 43876 40236 45052 40292
rect 45108 40236 45118 40292
rect 12684 40124 14252 40180
rect 14308 40124 14318 40180
rect 16818 40124 16828 40180
rect 16884 40124 18060 40180
rect 18116 40124 18126 40180
rect 18946 40124 18956 40180
rect 19012 40124 19292 40180
rect 19348 40124 19358 40180
rect 19506 40124 19516 40180
rect 19572 40124 19964 40180
rect 20020 40124 20030 40180
rect 20290 40124 20300 40180
rect 20356 40124 29260 40180
rect 29316 40124 29326 40180
rect 29586 40124 29596 40180
rect 29652 40124 29662 40180
rect 31042 40124 31052 40180
rect 31108 40124 31612 40180
rect 31668 40124 31678 40180
rect 31826 40124 31836 40180
rect 31892 40124 39228 40180
rect 39284 40124 39294 40180
rect 14466 40012 14476 40068
rect 14532 40012 18956 40068
rect 19012 40012 19022 40068
rect 19170 40012 19180 40068
rect 19236 40012 19516 40068
rect 19572 40012 19582 40068
rect 25778 40012 25788 40068
rect 25844 40012 30492 40068
rect 30548 40012 30558 40068
rect 40674 40012 40684 40068
rect 40740 40012 41244 40068
rect 41300 40012 41310 40068
rect 43138 40012 43148 40068
rect 43204 40012 43484 40068
rect 43540 40012 43550 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 19394 39900 19404 39956
rect 19460 39900 27356 39956
rect 27412 39900 27422 39956
rect 28578 39900 28588 39956
rect 28644 39900 30268 39956
rect 30324 39900 31612 39956
rect 31668 39900 31678 39956
rect 40786 39900 40796 39956
rect 40852 39900 41916 39956
rect 41972 39900 41982 39956
rect 16818 39788 16828 39844
rect 16884 39788 17164 39844
rect 17220 39788 20580 39844
rect 21634 39788 21644 39844
rect 21700 39788 23436 39844
rect 23492 39788 23502 39844
rect 25218 39788 25228 39844
rect 25284 39788 30828 39844
rect 30884 39788 30894 39844
rect 34178 39788 34188 39844
rect 34244 39788 35084 39844
rect 35140 39788 36876 39844
rect 36932 39788 36942 39844
rect 38434 39788 38444 39844
rect 38500 39788 43484 39844
rect 43540 39788 43550 39844
rect 20524 39732 20580 39788
rect 11554 39676 11564 39732
rect 11620 39676 14476 39732
rect 14532 39676 14542 39732
rect 19954 39676 19964 39732
rect 20020 39676 20188 39732
rect 20244 39676 20254 39732
rect 20524 39676 23884 39732
rect 23940 39676 24108 39732
rect 24164 39676 24174 39732
rect 28466 39676 28476 39732
rect 28532 39676 39116 39732
rect 39172 39676 39182 39732
rect 8754 39564 8764 39620
rect 8820 39564 9436 39620
rect 9492 39564 9502 39620
rect 12898 39564 12908 39620
rect 12964 39564 13580 39620
rect 13636 39564 13646 39620
rect 18386 39564 18396 39620
rect 18452 39564 20524 39620
rect 20580 39564 20590 39620
rect 21522 39564 21532 39620
rect 21588 39564 29372 39620
rect 29428 39564 29438 39620
rect 30258 39564 30268 39620
rect 30324 39564 30828 39620
rect 30884 39564 31388 39620
rect 31444 39564 31454 39620
rect 41794 39564 41804 39620
rect 41860 39564 42140 39620
rect 42196 39564 42206 39620
rect 43922 39564 43932 39620
rect 43988 39564 45388 39620
rect 45444 39564 46284 39620
rect 46340 39564 46620 39620
rect 46676 39564 46686 39620
rect 17602 39452 17612 39508
rect 17668 39452 18956 39508
rect 19012 39452 19022 39508
rect 24882 39452 24892 39508
rect 24948 39452 31164 39508
rect 31220 39452 31230 39508
rect 36418 39452 36428 39508
rect 36484 39452 37212 39508
rect 37268 39452 37278 39508
rect 37426 39452 37436 39508
rect 37492 39452 45164 39508
rect 45220 39452 45230 39508
rect 11442 39340 11452 39396
rect 11508 39340 12460 39396
rect 12516 39340 13804 39396
rect 13860 39340 13870 39396
rect 14354 39340 14364 39396
rect 14420 39340 20412 39396
rect 20468 39340 20478 39396
rect 23202 39340 23212 39396
rect 23268 39340 24220 39396
rect 24276 39340 24286 39396
rect 25106 39340 25116 39396
rect 25172 39340 25228 39396
rect 25284 39340 25294 39396
rect 29362 39340 29372 39396
rect 29428 39340 30380 39396
rect 30436 39340 31612 39396
rect 31668 39340 31678 39396
rect 39554 39340 39564 39396
rect 39620 39340 40572 39396
rect 40628 39340 41468 39396
rect 41524 39340 41534 39396
rect 42802 39340 42812 39396
rect 42868 39340 43820 39396
rect 43876 39340 43886 39396
rect 16818 39228 16828 39284
rect 16884 39228 18732 39284
rect 18788 39228 18798 39284
rect 19030 39228 19068 39284
rect 19124 39228 19134 39284
rect 20850 39228 20860 39284
rect 20916 39228 21756 39284
rect 21812 39228 31388 39284
rect 31444 39228 31454 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 11116 39116 11676 39172
rect 11732 39116 11742 39172
rect 20188 39116 23660 39172
rect 23716 39116 26236 39172
rect 26292 39116 26302 39172
rect 11116 38948 11172 39116
rect 20188 39060 20244 39116
rect 59200 39060 60000 39088
rect 11330 39004 11340 39060
rect 11396 39004 14028 39060
rect 14084 39004 14094 39060
rect 14802 39004 14812 39060
rect 14868 39004 16156 39060
rect 16212 39004 18284 39060
rect 18340 39004 18350 39060
rect 18498 39004 18508 39060
rect 18564 39004 20244 39060
rect 21074 39004 21084 39060
rect 21140 39004 21420 39060
rect 21476 39004 21486 39060
rect 22754 39004 22764 39060
rect 22820 39004 23996 39060
rect 24052 39004 26012 39060
rect 26068 39004 26078 39060
rect 26236 39004 26348 39060
rect 26404 39004 26414 39060
rect 29586 39004 29596 39060
rect 29652 39004 32956 39060
rect 33012 39004 33022 39060
rect 39778 39004 39788 39060
rect 39844 39004 41244 39060
rect 41300 39004 41310 39060
rect 46274 39004 46284 39060
rect 46340 39004 46732 39060
rect 46788 39004 46798 39060
rect 58258 39004 58268 39060
rect 58324 39004 60000 39060
rect 26236 38948 26292 39004
rect 59200 38976 60000 39004
rect 10882 38892 10892 38948
rect 10948 38892 13748 38948
rect 15138 38892 15148 38948
rect 15204 38892 16604 38948
rect 16660 38892 17276 38948
rect 17332 38892 24108 38948
rect 24164 38892 24174 38948
rect 26114 38892 26124 38948
rect 26180 38892 26292 38948
rect 26674 38892 26684 38948
rect 26740 38892 29148 38948
rect 29204 38892 29214 38948
rect 30594 38892 30604 38948
rect 30660 38892 30940 38948
rect 30996 38892 31006 38948
rect 43026 38892 43036 38948
rect 43092 38892 44044 38948
rect 44100 38892 44110 38948
rect 13692 38836 13748 38892
rect 10322 38780 10332 38836
rect 10388 38780 11452 38836
rect 11508 38780 11518 38836
rect 11778 38780 11788 38836
rect 11844 38780 13468 38836
rect 13524 38780 13534 38836
rect 13692 38780 16044 38836
rect 16100 38780 16110 38836
rect 18386 38780 18396 38836
rect 18452 38780 19628 38836
rect 19684 38780 23436 38836
rect 23492 38780 23502 38836
rect 23650 38780 23660 38836
rect 23716 38780 26572 38836
rect 26628 38780 26638 38836
rect 26852 38780 28140 38836
rect 28196 38780 28206 38836
rect 30818 38780 30828 38836
rect 30884 38780 31612 38836
rect 31668 38780 31678 38836
rect 41570 38780 41580 38836
rect 41636 38780 43596 38836
rect 43652 38780 44268 38836
rect 44324 38780 44334 38836
rect 46386 38780 46396 38836
rect 46452 38780 47404 38836
rect 47460 38780 47470 38836
rect 11452 38724 11508 38780
rect 26852 38724 26908 38780
rect 11452 38668 11900 38724
rect 11956 38668 11966 38724
rect 13234 38668 13244 38724
rect 13300 38668 20860 38724
rect 20916 38668 20926 38724
rect 24658 38668 24668 38724
rect 24724 38668 26124 38724
rect 26180 38668 26908 38724
rect 43250 38668 43260 38724
rect 43316 38668 46508 38724
rect 46564 38668 46574 38724
rect 20402 38556 20412 38612
rect 20468 38556 21308 38612
rect 21364 38556 21374 38612
rect 24434 38556 24444 38612
rect 24500 38556 25340 38612
rect 25396 38556 25406 38612
rect 33394 38556 33404 38612
rect 33460 38556 37996 38612
rect 38052 38556 38062 38612
rect 42130 38556 42140 38612
rect 42196 38556 43932 38612
rect 43988 38556 43998 38612
rect 26898 38444 26908 38500
rect 26964 38444 27804 38500
rect 27860 38444 27870 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 59200 38388 60000 38416
rect 14690 38332 14700 38388
rect 14756 38332 24332 38388
rect 24388 38332 24398 38388
rect 25666 38332 25676 38388
rect 25732 38332 26348 38388
rect 26404 38332 26414 38388
rect 58146 38332 58156 38388
rect 58212 38332 60000 38388
rect 59200 38304 60000 38332
rect 15894 38220 15932 38276
rect 15988 38220 15998 38276
rect 20962 38220 20972 38276
rect 21028 38220 31500 38276
rect 31556 38220 32844 38276
rect 32900 38220 32910 38276
rect 12898 38108 12908 38164
rect 12964 38108 13916 38164
rect 13972 38108 13982 38164
rect 15698 38108 15708 38164
rect 15764 38108 19292 38164
rect 19348 38108 19740 38164
rect 19796 38108 19806 38164
rect 22866 38108 22876 38164
rect 22932 38108 23324 38164
rect 23380 38108 24108 38164
rect 24164 38108 24444 38164
rect 24500 38108 24510 38164
rect 24994 38108 25004 38164
rect 25060 38108 31612 38164
rect 31668 38108 31948 38164
rect 32274 38108 32284 38164
rect 32340 38108 34300 38164
rect 34356 38108 34412 38164
rect 34468 38108 34478 38164
rect 31892 38052 31948 38108
rect 13794 37996 13804 38052
rect 13860 37996 14028 38052
rect 14084 37996 15148 38052
rect 16034 37996 16044 38052
rect 16100 37996 16492 38052
rect 16548 37996 16558 38052
rect 17154 37996 17164 38052
rect 17220 37996 17230 38052
rect 19618 37996 19628 38052
rect 19684 37996 22764 38052
rect 22820 37996 22830 38052
rect 23202 37996 23212 38052
rect 23268 37996 24892 38052
rect 24948 37996 24958 38052
rect 25330 37996 25340 38052
rect 25396 37996 26012 38052
rect 26068 37996 26078 38052
rect 31892 37996 32620 38052
rect 32676 37996 32686 38052
rect 34514 37996 34524 38052
rect 34580 37996 35084 38052
rect 35140 37996 35150 38052
rect 49522 37996 49532 38052
rect 49588 37996 55580 38052
rect 55636 37996 55646 38052
rect 15092 37940 15148 37996
rect 17164 37940 17220 37996
rect 9650 37884 9660 37940
rect 9716 37884 10444 37940
rect 10500 37884 11116 37940
rect 11172 37884 11182 37940
rect 15092 37884 17220 37940
rect 19730 37884 19740 37940
rect 19796 37884 23828 37940
rect 24098 37884 24108 37940
rect 24164 37884 25900 37940
rect 25956 37884 25966 37940
rect 27906 37884 27916 37940
rect 27972 37884 29260 37940
rect 29316 37884 29326 37940
rect 31938 37884 31948 37940
rect 32004 37884 33964 37940
rect 34020 37884 34030 37940
rect 34626 37884 34636 37940
rect 34692 37884 42476 37940
rect 42532 37884 42542 37940
rect 23772 37828 23828 37884
rect 1698 37772 1708 37828
rect 1764 37772 1774 37828
rect 11732 37772 19404 37828
rect 19460 37772 19470 37828
rect 21970 37772 21980 37828
rect 22036 37772 23548 37828
rect 23604 37772 23614 37828
rect 23772 37772 24332 37828
rect 24388 37772 24398 37828
rect 24658 37772 24668 37828
rect 24724 37772 32732 37828
rect 32788 37772 32798 37828
rect 35634 37772 35644 37828
rect 35700 37772 37212 37828
rect 37268 37772 37278 37828
rect 0 37716 800 37744
rect 1708 37716 1764 37772
rect 0 37660 1764 37716
rect 0 37632 800 37660
rect 11732 37604 11788 37772
rect 59200 37716 60000 37744
rect 18050 37660 18060 37716
rect 18116 37660 18508 37716
rect 18564 37660 18574 37716
rect 22754 37660 22764 37716
rect 22820 37660 24780 37716
rect 24836 37660 24846 37716
rect 25106 37660 25116 37716
rect 25172 37660 25956 37716
rect 26338 37660 26348 37716
rect 26404 37660 26684 37716
rect 26740 37660 26750 37716
rect 29362 37660 29372 37716
rect 29428 37660 30716 37716
rect 30772 37660 30782 37716
rect 57922 37660 57932 37716
rect 57988 37660 60000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 25900 37604 25956 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37632 60000 37660
rect 8978 37548 8988 37604
rect 9044 37548 11788 37604
rect 15092 37548 18620 37604
rect 18676 37548 18686 37604
rect 18834 37548 18844 37604
rect 18900 37548 19572 37604
rect 20402 37548 20412 37604
rect 20468 37548 21980 37604
rect 22036 37548 22046 37604
rect 24322 37548 24332 37604
rect 24388 37548 25116 37604
rect 25172 37548 25182 37604
rect 25900 37548 28252 37604
rect 28308 37548 28318 37604
rect 34290 37548 34300 37604
rect 34356 37548 36988 37604
rect 37044 37548 37054 37604
rect 15092 37492 15148 37548
rect 19516 37492 19572 37548
rect 12114 37436 12124 37492
rect 12180 37436 15148 37492
rect 15810 37436 15820 37492
rect 15876 37436 18620 37492
rect 18676 37436 18956 37492
rect 19012 37436 19022 37492
rect 19506 37436 19516 37492
rect 19572 37436 23772 37492
rect 23828 37436 25564 37492
rect 25620 37436 25630 37492
rect 41906 37436 41916 37492
rect 41972 37436 45836 37492
rect 45892 37436 46844 37492
rect 46900 37436 46910 37492
rect 14214 37324 14252 37380
rect 14308 37324 26796 37380
rect 26852 37324 27468 37380
rect 27524 37324 27534 37380
rect 38546 37324 38556 37380
rect 38612 37324 39340 37380
rect 39396 37324 39788 37380
rect 39844 37324 39854 37380
rect 7858 37212 7868 37268
rect 7924 37212 10556 37268
rect 10612 37212 10892 37268
rect 10948 37212 10958 37268
rect 12786 37212 12796 37268
rect 12852 37212 15820 37268
rect 15876 37212 15886 37268
rect 16034 37212 16044 37268
rect 16100 37212 19292 37268
rect 19348 37212 19358 37268
rect 19506 37212 19516 37268
rect 19572 37212 20412 37268
rect 20468 37212 20478 37268
rect 24322 37212 24332 37268
rect 24388 37212 26908 37268
rect 26964 37212 26974 37268
rect 33170 37212 33180 37268
rect 33236 37212 34412 37268
rect 34468 37212 35196 37268
rect 35252 37212 35262 37268
rect 39554 37212 39564 37268
rect 39620 37212 40908 37268
rect 40964 37212 40974 37268
rect 9650 37100 9660 37156
rect 9716 37100 11228 37156
rect 11284 37100 11294 37156
rect 16044 37044 16100 37212
rect 17490 37100 17500 37156
rect 17556 37100 19852 37156
rect 19908 37100 19918 37156
rect 21746 37100 21756 37156
rect 21812 37100 22820 37156
rect 30230 37100 30268 37156
rect 30324 37100 30716 37156
rect 30772 37100 31612 37156
rect 31668 37100 32396 37156
rect 32452 37100 32462 37156
rect 34178 37100 34188 37156
rect 34244 37100 34748 37156
rect 34804 37100 35420 37156
rect 35476 37100 35756 37156
rect 35812 37100 35822 37156
rect 40002 37100 40012 37156
rect 40068 37100 41804 37156
rect 41860 37100 41870 37156
rect 22764 37044 22820 37100
rect 12898 36988 12908 37044
rect 12964 36988 16100 37044
rect 17714 36988 17724 37044
rect 17780 36988 18844 37044
rect 18900 36988 18910 37044
rect 19618 36988 19628 37044
rect 19684 36988 20300 37044
rect 20356 36988 20366 37044
rect 20514 36988 20524 37044
rect 20580 36988 21980 37044
rect 22036 36988 22046 37044
rect 22754 36988 22764 37044
rect 22820 36988 29820 37044
rect 29876 36988 29886 37044
rect 33730 36988 33740 37044
rect 33796 36988 34972 37044
rect 35028 36988 35038 37044
rect 39890 36988 39900 37044
rect 39956 36988 41132 37044
rect 41188 36988 41198 37044
rect 10098 36876 10108 36932
rect 10164 36876 11452 36932
rect 11508 36876 11518 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 18396 36820 18452 36988
rect 24434 36876 24444 36932
rect 24500 36876 25564 36932
rect 25620 36876 25630 36932
rect 27346 36876 27356 36932
rect 27412 36876 27468 36932
rect 27524 36876 27534 36932
rect 28354 36876 28364 36932
rect 28420 36876 31052 36932
rect 31108 36876 31500 36932
rect 31556 36876 31566 36932
rect 36866 36876 36876 36932
rect 36932 36876 42812 36932
rect 42868 36876 42878 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 18386 36764 18396 36820
rect 18452 36764 18462 36820
rect 18946 36764 18956 36820
rect 19012 36764 32172 36820
rect 32228 36764 32238 36820
rect 17602 36652 17612 36708
rect 17668 36652 21868 36708
rect 21924 36652 21934 36708
rect 25106 36652 25116 36708
rect 25172 36652 33516 36708
rect 33572 36652 33582 36708
rect 37874 36652 37884 36708
rect 37940 36652 40012 36708
rect 40068 36652 40078 36708
rect 18610 36540 18620 36596
rect 18676 36540 18844 36596
rect 18900 36540 18910 36596
rect 24444 36540 25340 36596
rect 25396 36540 25406 36596
rect 26012 36540 26572 36596
rect 26628 36540 29260 36596
rect 29316 36540 29326 36596
rect 43810 36540 43820 36596
rect 43876 36540 45612 36596
rect 45668 36540 47068 36596
rect 47124 36540 47134 36596
rect 24444 36484 24500 36540
rect 26012 36484 26068 36540
rect 12450 36428 12460 36484
rect 12516 36428 14140 36484
rect 14196 36428 15820 36484
rect 15876 36428 16716 36484
rect 16772 36428 16782 36484
rect 18610 36428 18620 36484
rect 18676 36428 19404 36484
rect 19460 36428 19470 36484
rect 19852 36428 20188 36484
rect 20244 36428 20254 36484
rect 21746 36428 21756 36484
rect 21812 36428 23548 36484
rect 23604 36428 23614 36484
rect 24434 36428 24444 36484
rect 24500 36428 24510 36484
rect 26002 36428 26012 36484
rect 26068 36428 26078 36484
rect 27906 36428 27916 36484
rect 27972 36428 30156 36484
rect 30212 36428 30222 36484
rect 30930 36428 30940 36484
rect 30996 36428 33068 36484
rect 33124 36428 33134 36484
rect 34626 36428 34636 36484
rect 34692 36428 35644 36484
rect 35700 36428 35710 36484
rect 36866 36428 36876 36484
rect 36932 36428 37884 36484
rect 37940 36428 37950 36484
rect 39106 36428 39116 36484
rect 39172 36428 40124 36484
rect 40180 36428 40908 36484
rect 40964 36428 40974 36484
rect 42802 36428 42812 36484
rect 42868 36428 44044 36484
rect 44100 36428 44110 36484
rect 19852 36372 19908 36428
rect 59200 36372 60000 36400
rect 9314 36316 9324 36372
rect 9380 36316 9996 36372
rect 10052 36316 10062 36372
rect 10994 36316 11004 36372
rect 11060 36316 12572 36372
rect 12628 36316 12638 36372
rect 13234 36316 13244 36372
rect 13300 36316 19908 36372
rect 20066 36316 20076 36372
rect 20132 36316 24556 36372
rect 24612 36316 24622 36372
rect 26348 36316 32508 36372
rect 32564 36316 32574 36372
rect 35522 36316 35532 36372
rect 35588 36316 37996 36372
rect 38052 36316 38062 36372
rect 41570 36316 41580 36372
rect 41636 36316 45836 36372
rect 45892 36316 46844 36372
rect 46900 36316 46910 36372
rect 57810 36316 57820 36372
rect 57876 36316 60000 36372
rect 11004 36260 11060 36316
rect 26348 36260 26404 36316
rect 59200 36288 60000 36316
rect 9202 36204 9212 36260
rect 9268 36204 11060 36260
rect 11442 36204 11452 36260
rect 11508 36204 11518 36260
rect 19282 36204 19292 36260
rect 19348 36204 26404 36260
rect 26786 36204 26796 36260
rect 26852 36204 27580 36260
rect 27636 36204 27646 36260
rect 30594 36204 30604 36260
rect 30660 36204 30940 36260
rect 30996 36204 31006 36260
rect 43026 36204 43036 36260
rect 43092 36204 44156 36260
rect 44212 36204 44222 36260
rect 11452 36148 11508 36204
rect 26796 36148 26852 36204
rect 11452 36092 15708 36148
rect 15764 36092 16100 36148
rect 17378 36092 17388 36148
rect 17444 36092 19628 36148
rect 19684 36092 19694 36148
rect 20178 36092 20188 36148
rect 20244 36092 26852 36148
rect 37986 36092 37996 36148
rect 38052 36092 38892 36148
rect 38948 36092 38958 36148
rect 16044 35924 16100 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 20962 35980 20972 36036
rect 21028 35980 23660 36036
rect 23716 35980 24220 36036
rect 24276 35980 24286 36036
rect 25078 35980 25116 36036
rect 25172 35980 25182 36036
rect 30258 35980 30268 36036
rect 30324 35980 30940 36036
rect 30996 35980 32060 36036
rect 32116 35980 32126 36036
rect 34178 35980 34188 36036
rect 34244 35980 41916 36036
rect 41972 35980 43708 36036
rect 43764 35980 43774 36036
rect 14578 35868 14588 35924
rect 14644 35868 15148 35924
rect 16044 35868 20300 35924
rect 20356 35868 20366 35924
rect 23538 35868 23548 35924
rect 23604 35868 24444 35924
rect 24500 35868 24510 35924
rect 26562 35868 26572 35924
rect 26628 35868 27020 35924
rect 27076 35868 27086 35924
rect 29026 35868 29036 35924
rect 29092 35868 33852 35924
rect 33908 35868 34524 35924
rect 34580 35868 34590 35924
rect 34850 35868 34860 35924
rect 34916 35868 35644 35924
rect 35700 35868 36204 35924
rect 36260 35868 36270 35924
rect 38770 35868 38780 35924
rect 38836 35868 39676 35924
rect 39732 35868 42028 35924
rect 42084 35868 42094 35924
rect 8306 35756 8316 35812
rect 8372 35756 9548 35812
rect 9604 35756 10724 35812
rect 11330 35756 11340 35812
rect 11396 35756 11676 35812
rect 11732 35756 12348 35812
rect 12404 35756 13692 35812
rect 13748 35756 13758 35812
rect 10668 35588 10724 35756
rect 15092 35700 15148 35868
rect 28924 35756 31724 35812
rect 31780 35756 31790 35812
rect 31892 35756 34972 35812
rect 35028 35756 36428 35812
rect 36484 35756 36494 35812
rect 46722 35756 46732 35812
rect 46788 35756 55580 35812
rect 55636 35756 55646 35812
rect 28924 35700 28980 35756
rect 31892 35700 31948 35756
rect 59200 35700 60000 35728
rect 10882 35644 10892 35700
rect 10948 35644 11900 35700
rect 11956 35644 11966 35700
rect 15092 35644 18508 35700
rect 18564 35644 18574 35700
rect 23426 35644 23436 35700
rect 23492 35644 25340 35700
rect 25396 35644 25406 35700
rect 27346 35644 27356 35700
rect 27412 35644 28924 35700
rect 28980 35644 28990 35700
rect 31378 35644 31388 35700
rect 31444 35644 31948 35700
rect 57922 35644 57932 35700
rect 57988 35644 60000 35700
rect 59200 35616 60000 35644
rect 10668 35532 11788 35588
rect 11844 35532 14028 35588
rect 14084 35532 14588 35588
rect 14644 35532 14654 35588
rect 18050 35532 18060 35588
rect 18116 35532 21420 35588
rect 21476 35532 21486 35588
rect 24098 35532 24108 35588
rect 24164 35532 24668 35588
rect 24724 35532 24734 35588
rect 29810 35532 29820 35588
rect 29876 35532 30604 35588
rect 30660 35532 30670 35588
rect 16594 35420 16604 35476
rect 16660 35420 17836 35476
rect 17892 35420 19292 35476
rect 19348 35420 21868 35476
rect 21924 35420 21934 35476
rect 30034 35420 30044 35476
rect 30100 35420 33628 35476
rect 33684 35420 34636 35476
rect 34692 35420 34702 35476
rect 18022 35308 18060 35364
rect 18116 35308 18126 35364
rect 23548 35308 25564 35364
rect 25620 35308 25630 35364
rect 26674 35308 26684 35364
rect 26740 35308 28364 35364
rect 28420 35308 29260 35364
rect 29316 35308 29326 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 23548 35252 23604 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 12898 35196 12908 35252
rect 12964 35196 13468 35252
rect 13524 35196 14700 35252
rect 14756 35196 14766 35252
rect 19170 35196 19180 35252
rect 19236 35196 23604 35252
rect 26226 35196 26236 35252
rect 26292 35196 31276 35252
rect 31332 35196 32732 35252
rect 32788 35196 32798 35252
rect 27458 35084 27468 35140
rect 27524 35084 28476 35140
rect 28532 35084 28542 35140
rect 31378 35084 31388 35140
rect 31444 35084 31948 35140
rect 34962 35084 34972 35140
rect 35028 35084 35980 35140
rect 36036 35084 36046 35140
rect 8372 34972 10780 35028
rect 10836 34972 10846 35028
rect 11554 34972 11564 35028
rect 11620 34972 19964 35028
rect 20020 34972 20636 35028
rect 20692 34972 20702 35028
rect 22530 34972 22540 35028
rect 22596 34972 28140 35028
rect 28196 34972 29260 35028
rect 29316 34972 29326 35028
rect 31892 34972 31948 35084
rect 32004 34972 32396 35028
rect 32452 34972 32462 35028
rect 40002 34972 40012 35028
rect 40068 34972 44156 35028
rect 44212 34972 44222 35028
rect 8372 34692 8428 34972
rect 8978 34860 8988 34916
rect 9044 34860 9996 34916
rect 10052 34860 10062 34916
rect 14914 34860 14924 34916
rect 14980 34860 16044 34916
rect 16100 34860 16110 34916
rect 22194 34860 22204 34916
rect 22260 34860 23436 34916
rect 23492 34860 23502 34916
rect 25778 34860 25788 34916
rect 25844 34860 26684 34916
rect 26740 34860 29148 34916
rect 29204 34860 29484 34916
rect 29540 34860 31164 34916
rect 31220 34860 31230 34916
rect 35074 34860 35084 34916
rect 35140 34860 35868 34916
rect 35924 34860 35934 34916
rect 45378 34860 45388 34916
rect 45444 34860 55580 34916
rect 55636 34860 55646 34916
rect 12226 34748 12236 34804
rect 12292 34748 12908 34804
rect 12964 34748 15036 34804
rect 15092 34748 16492 34804
rect 16548 34748 16558 34804
rect 18610 34748 18620 34804
rect 18676 34748 19180 34804
rect 19236 34748 19404 34804
rect 19460 34748 19470 34804
rect 28466 34748 28476 34804
rect 28532 34748 30380 34804
rect 30436 34748 30446 34804
rect 32498 34748 32508 34804
rect 32564 34748 40012 34804
rect 40068 34748 40078 34804
rect 8082 34636 8092 34692
rect 8148 34636 8428 34692
rect 12562 34636 12572 34692
rect 12628 34636 13580 34692
rect 13636 34636 13646 34692
rect 16818 34636 16828 34692
rect 16884 34636 17948 34692
rect 18004 34636 18014 34692
rect 25442 34636 25452 34692
rect 25508 34636 27020 34692
rect 27076 34636 27086 34692
rect 34626 34636 34636 34692
rect 34692 34636 34860 34692
rect 34916 34636 34926 34692
rect 24658 34524 24668 34580
rect 24724 34524 25900 34580
rect 25956 34524 30716 34580
rect 30772 34524 31164 34580
rect 31220 34524 31230 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 20290 34412 20300 34468
rect 20356 34412 25788 34468
rect 25844 34412 26684 34468
rect 26740 34412 26750 34468
rect 15698 34300 15708 34356
rect 15764 34300 17724 34356
rect 17780 34300 18844 34356
rect 18900 34300 18910 34356
rect 33394 34300 33404 34356
rect 33460 34300 33852 34356
rect 33908 34300 38108 34356
rect 38164 34300 38174 34356
rect 8530 34188 8540 34244
rect 8596 34188 10444 34244
rect 10500 34188 10668 34244
rect 10724 34188 10734 34244
rect 16482 34188 16492 34244
rect 16548 34188 19852 34244
rect 19908 34188 19918 34244
rect 22306 34188 22316 34244
rect 22372 34188 23772 34244
rect 23828 34188 24444 34244
rect 24500 34188 26012 34244
rect 26068 34188 26078 34244
rect 4162 34076 4172 34132
rect 4228 34076 4844 34132
rect 4900 34076 4910 34132
rect 10882 34076 10892 34132
rect 10948 34076 13580 34132
rect 13636 34076 13646 34132
rect 20626 34076 20636 34132
rect 20692 34076 22652 34132
rect 22708 34076 22718 34132
rect 24770 34076 24780 34132
rect 24836 34076 25452 34132
rect 25508 34076 25518 34132
rect 26338 34076 26348 34132
rect 26404 34076 29036 34132
rect 29092 34076 29102 34132
rect 32162 34076 32172 34132
rect 32228 34076 34412 34132
rect 34468 34076 34478 34132
rect 36978 34076 36988 34132
rect 37044 34076 39116 34132
rect 39172 34076 39182 34132
rect 39778 34076 39788 34132
rect 39844 34076 40348 34132
rect 40404 34076 41132 34132
rect 41188 34076 41198 34132
rect 44146 34076 44156 34132
rect 44212 34076 45388 34132
rect 45444 34076 45454 34132
rect 34412 34020 34468 34076
rect 20962 33964 20972 34020
rect 21028 33964 26124 34020
rect 26180 33964 26190 34020
rect 26348 33964 29820 34020
rect 29876 33964 30716 34020
rect 30772 33964 30782 34020
rect 34412 33964 38668 34020
rect 38724 33964 40908 34020
rect 40964 33964 40974 34020
rect 43474 33964 43484 34020
rect 43540 33964 44604 34020
rect 44660 33964 45276 34020
rect 45332 33964 45342 34020
rect 26348 33908 26404 33964
rect 1922 33852 1932 33908
rect 1988 33852 1998 33908
rect 14578 33852 14588 33908
rect 14644 33852 15372 33908
rect 15428 33852 15438 33908
rect 23202 33852 23212 33908
rect 23268 33852 26404 33908
rect 26674 33852 26684 33908
rect 26740 33852 28700 33908
rect 28756 33852 28766 33908
rect 0 33684 800 33712
rect 1932 33684 1988 33852
rect 13682 33740 13692 33796
rect 13748 33740 22876 33796
rect 22932 33740 22942 33796
rect 24882 33740 24892 33796
rect 24948 33740 25676 33796
rect 25732 33740 25742 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 59200 33684 60000 33712
rect 0 33628 1988 33684
rect 4834 33628 4844 33684
rect 4900 33628 5796 33684
rect 11666 33628 11676 33684
rect 11732 33628 21756 33684
rect 21812 33628 22316 33684
rect 22372 33628 22382 33684
rect 23426 33628 23436 33684
rect 23492 33628 27132 33684
rect 27188 33628 27198 33684
rect 58146 33628 58156 33684
rect 58212 33628 60000 33684
rect 0 33600 800 33628
rect 5740 33572 5796 33628
rect 59200 33600 60000 33628
rect 5740 33516 18564 33572
rect 18834 33516 18844 33572
rect 18900 33516 19516 33572
rect 19572 33516 19582 33572
rect 20290 33516 20300 33572
rect 20356 33516 21308 33572
rect 21364 33516 21374 33572
rect 23874 33516 23884 33572
rect 23940 33516 24668 33572
rect 24724 33516 25676 33572
rect 25732 33516 25742 33572
rect 18508 33460 18564 33516
rect 14466 33404 14476 33460
rect 14532 33404 16660 33460
rect 18508 33404 24500 33460
rect 25330 33404 25340 33460
rect 25396 33404 28140 33460
rect 28196 33404 28364 33460
rect 28420 33404 28430 33460
rect 35644 33404 38220 33460
rect 38276 33404 38286 33460
rect 16604 33348 16660 33404
rect 4274 33292 4284 33348
rect 4340 33292 8876 33348
rect 8932 33292 8942 33348
rect 9986 33292 9996 33348
rect 10052 33292 10780 33348
rect 10836 33292 10846 33348
rect 12674 33292 12684 33348
rect 12740 33292 16436 33348
rect 16594 33292 16604 33348
rect 16660 33292 20300 33348
rect 20356 33292 20366 33348
rect 20738 33292 20748 33348
rect 20804 33292 21756 33348
rect 21812 33292 22652 33348
rect 22708 33292 23100 33348
rect 23156 33292 23324 33348
rect 23380 33292 23390 33348
rect 24210 33292 24220 33348
rect 24276 33292 24286 33348
rect 16380 33236 16436 33292
rect 10546 33180 10556 33236
rect 10612 33180 14252 33236
rect 14308 33180 14700 33236
rect 14756 33180 14766 33236
rect 15092 33180 15596 33236
rect 15652 33180 15662 33236
rect 16380 33180 17052 33236
rect 17108 33180 17118 33236
rect 18610 33180 18620 33236
rect 18676 33180 19180 33236
rect 19236 33180 20188 33236
rect 20244 33180 20254 33236
rect 15092 33124 15148 33180
rect 24220 33124 24276 33292
rect 24444 33236 24500 33404
rect 35644 33348 35700 33404
rect 30370 33292 30380 33348
rect 30436 33292 30940 33348
rect 30996 33292 31006 33348
rect 32162 33292 32172 33348
rect 32228 33292 33068 33348
rect 33124 33292 35644 33348
rect 35700 33292 35710 33348
rect 37314 33292 37324 33348
rect 37380 33292 45052 33348
rect 45108 33292 45118 33348
rect 24444 33180 27580 33236
rect 27636 33180 28476 33236
rect 28532 33180 28542 33236
rect 40338 33180 40348 33236
rect 40404 33180 41356 33236
rect 41412 33180 42140 33236
rect 42196 33180 42206 33236
rect 12114 33068 12124 33124
rect 12180 33068 13356 33124
rect 13412 33068 15148 33124
rect 18498 33068 18508 33124
rect 18564 33068 19292 33124
rect 19348 33068 19358 33124
rect 20738 33068 20748 33124
rect 20804 33068 22204 33124
rect 22260 33068 23324 33124
rect 23380 33068 23660 33124
rect 23716 33068 23726 33124
rect 24220 33068 26908 33124
rect 26964 33068 29708 33124
rect 29764 33068 29774 33124
rect 0 33012 800 33040
rect 59200 33012 60000 33040
rect 0 32956 1932 33012
rect 1988 32956 1998 33012
rect 16594 32956 16604 33012
rect 16660 32956 18844 33012
rect 18900 32956 19684 33012
rect 23202 32956 23212 33012
rect 23268 32956 28140 33012
rect 28196 32956 28206 33012
rect 58146 32956 58156 33012
rect 58212 32956 60000 33012
rect 0 32928 800 32956
rect 11218 32844 11228 32900
rect 11284 32844 15372 32900
rect 15428 32844 17836 32900
rect 17892 32844 17902 32900
rect 19366 32844 19404 32900
rect 19460 32844 19470 32900
rect 19628 32788 19684 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 59200 32928 60000 32956
rect 22204 32844 25228 32900
rect 25284 32844 26572 32900
rect 26628 32844 26638 32900
rect 15922 32732 15932 32788
rect 15988 32732 17948 32788
rect 18004 32732 18014 32788
rect 18946 32732 18956 32788
rect 19012 32732 19292 32788
rect 19348 32732 19358 32788
rect 19628 32732 21532 32788
rect 21588 32732 21598 32788
rect 22204 32676 22260 32844
rect 22418 32732 22428 32788
rect 22484 32732 24108 32788
rect 24164 32732 25452 32788
rect 25508 32732 25518 32788
rect 30342 32732 30380 32788
rect 30436 32732 30446 32788
rect 37212 32732 38668 32788
rect 38724 32732 39004 32788
rect 39060 32732 39070 32788
rect 37212 32676 37268 32732
rect 13570 32620 13580 32676
rect 13636 32620 15148 32676
rect 15204 32620 15708 32676
rect 15764 32620 15774 32676
rect 16482 32620 16492 32676
rect 16548 32620 22260 32676
rect 22866 32620 22876 32676
rect 22932 32620 24668 32676
rect 24724 32620 24734 32676
rect 31602 32620 31612 32676
rect 31668 32620 36876 32676
rect 36932 32620 37212 32676
rect 37268 32620 37278 32676
rect 38322 32620 38332 32676
rect 38388 32620 39732 32676
rect 39676 32564 39732 32620
rect 8866 32508 8876 32564
rect 8932 32508 10220 32564
rect 10276 32508 10668 32564
rect 10724 32508 11788 32564
rect 11844 32508 11854 32564
rect 12450 32508 12460 32564
rect 12516 32508 14028 32564
rect 14084 32508 14588 32564
rect 14644 32508 14654 32564
rect 17042 32508 17052 32564
rect 17108 32508 19964 32564
rect 20020 32508 21308 32564
rect 21364 32508 21374 32564
rect 38210 32508 38220 32564
rect 38276 32508 39228 32564
rect 39284 32508 39294 32564
rect 39666 32508 39676 32564
rect 39732 32508 39742 32564
rect 13458 32396 13468 32452
rect 13524 32396 14140 32452
rect 14196 32396 14206 32452
rect 15138 32396 15148 32452
rect 15204 32396 24108 32452
rect 24164 32396 24174 32452
rect 37874 32396 37884 32452
rect 37940 32396 38892 32452
rect 38948 32396 38958 32452
rect 0 32340 800 32368
rect 0 32284 1708 32340
rect 1764 32284 1774 32340
rect 0 32256 800 32284
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 11106 32060 11116 32116
rect 11172 32060 21756 32116
rect 21812 32060 21822 32116
rect 12786 31948 12796 32004
rect 12852 31948 14308 32004
rect 14252 31892 14308 31948
rect 1922 31836 1932 31892
rect 1988 31836 1998 31892
rect 10546 31836 10556 31892
rect 10612 31836 14308 31892
rect 14690 31836 14700 31892
rect 14756 31836 17164 31892
rect 17220 31836 17230 31892
rect 18274 31836 18284 31892
rect 18340 31836 18844 31892
rect 18900 31836 19068 31892
rect 19124 31836 19134 31892
rect 23958 31836 23996 31892
rect 24052 31836 24062 31892
rect 0 31668 800 31696
rect 1932 31668 1988 31836
rect 8978 31724 8988 31780
rect 9044 31724 9996 31780
rect 10052 31724 10892 31780
rect 10948 31724 10958 31780
rect 19282 31724 19292 31780
rect 19348 31724 28028 31780
rect 28084 31724 28094 31780
rect 0 31612 1988 31668
rect 8754 31612 8764 31668
rect 8820 31612 14700 31668
rect 14756 31612 15596 31668
rect 15652 31612 15662 31668
rect 23650 31612 23660 31668
rect 23716 31612 25452 31668
rect 25508 31612 25518 31668
rect 26852 31612 29596 31668
rect 29652 31612 29662 31668
rect 0 31584 800 31612
rect 14354 31500 14364 31556
rect 14420 31500 23548 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 23492 31332 23548 31500
rect 26852 31444 26908 31612
rect 24770 31388 24780 31444
rect 24836 31388 25116 31444
rect 25172 31388 26908 31444
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 16370 31276 16380 31332
rect 16436 31276 19460 31332
rect 23492 31276 30268 31332
rect 30324 31276 30334 31332
rect 19404 31220 19460 31276
rect 9874 31164 9884 31220
rect 9940 31164 12348 31220
rect 12404 31164 15820 31220
rect 15876 31164 15886 31220
rect 16706 31164 16716 31220
rect 16772 31164 19180 31220
rect 19236 31164 19246 31220
rect 19404 31164 19740 31220
rect 19796 31164 20300 31220
rect 20356 31164 20366 31220
rect 23426 31164 23436 31220
rect 23492 31164 24444 31220
rect 24500 31164 24892 31220
rect 24948 31164 24958 31220
rect 8530 31052 8540 31108
rect 8596 31052 9548 31108
rect 9604 31052 9614 31108
rect 18050 31052 18060 31108
rect 18116 31052 19628 31108
rect 19684 31052 19694 31108
rect 41906 31052 41916 31108
rect 41972 31052 57820 31108
rect 57876 31052 57886 31108
rect 0 30996 800 31024
rect 0 30940 1988 30996
rect 6066 30940 6076 30996
rect 6132 30940 18172 30996
rect 18228 30940 18238 30996
rect 30146 30940 30156 30996
rect 30212 30940 31500 30996
rect 31556 30940 32956 30996
rect 33012 30940 33022 30996
rect 0 30912 800 30940
rect 1932 30884 1988 30940
rect 1922 30828 1932 30884
rect 1988 30828 1998 30884
rect 20962 30828 20972 30884
rect 21028 30828 21756 30884
rect 21812 30828 22316 30884
rect 22372 30828 22764 30884
rect 22820 30828 22830 30884
rect 24658 30828 24668 30884
rect 24724 30828 25340 30884
rect 25396 30828 25406 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 4274 30380 4284 30436
rect 4340 30380 9100 30436
rect 9156 30380 12572 30436
rect 12628 30380 12638 30436
rect 14578 30380 14588 30436
rect 14644 30380 33068 30436
rect 33124 30380 33134 30436
rect 0 30324 800 30352
rect 59200 30324 60000 30352
rect 0 30268 1708 30324
rect 1764 30268 1774 30324
rect 17378 30268 17388 30324
rect 17444 30268 17948 30324
rect 18004 30268 18014 30324
rect 24322 30268 24332 30324
rect 24388 30268 25116 30324
rect 25172 30268 25182 30324
rect 36194 30268 36204 30324
rect 36260 30268 36988 30324
rect 37044 30268 37054 30324
rect 58146 30268 58156 30324
rect 58212 30268 60000 30324
rect 0 30240 800 30268
rect 59200 30240 60000 30268
rect 12226 30156 12236 30212
rect 12292 30156 17836 30212
rect 17892 30156 17902 30212
rect 19628 30156 24556 30212
rect 24612 30156 25452 30212
rect 25508 30156 26908 30212
rect 34290 30156 34300 30212
rect 34356 30156 34748 30212
rect 34804 30156 35532 30212
rect 35588 30156 35598 30212
rect 19628 30100 19684 30156
rect 26852 30100 26908 30156
rect 18274 30044 18284 30100
rect 18340 30044 18732 30100
rect 18788 30044 18798 30100
rect 18946 30044 18956 30100
rect 19012 30044 19628 30100
rect 19684 30044 19694 30100
rect 20402 30044 20412 30100
rect 20468 30044 22988 30100
rect 23044 30044 23054 30100
rect 23650 30044 23660 30100
rect 23716 30044 25004 30100
rect 25060 30044 25788 30100
rect 25844 30044 25854 30100
rect 26852 30044 31612 30100
rect 31668 30044 31678 30100
rect 34850 30044 34860 30100
rect 34916 30044 41916 30100
rect 41972 30044 41982 30100
rect 15250 29932 15260 29988
rect 15316 29932 16492 29988
rect 16548 29932 16558 29988
rect 19058 29932 19068 29988
rect 19124 29932 20972 29988
rect 21028 29932 21038 29988
rect 24434 29932 24444 29988
rect 24500 29932 25116 29988
rect 25172 29932 26684 29988
rect 26740 29932 26750 29988
rect 0 29652 800 29680
rect 0 29596 2156 29652
rect 2212 29596 2222 29652
rect 8306 29596 8316 29652
rect 8372 29596 11788 29652
rect 11844 29596 12348 29652
rect 12404 29596 12414 29652
rect 0 29568 800 29596
rect 15260 29540 15316 29932
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 35858 29708 35868 29764
rect 35924 29708 36876 29764
rect 36932 29708 38108 29764
rect 38164 29708 38174 29764
rect 28578 29596 28588 29652
rect 28644 29596 34412 29652
rect 34468 29596 34478 29652
rect 4274 29484 4284 29540
rect 4340 29484 15316 29540
rect 10098 29372 10108 29428
rect 10164 29372 16772 29428
rect 20626 29372 20636 29428
rect 20692 29372 22092 29428
rect 22148 29372 22158 29428
rect 31266 29372 31276 29428
rect 31332 29372 33628 29428
rect 33684 29372 33694 29428
rect 38882 29372 38892 29428
rect 38948 29372 41580 29428
rect 41636 29372 41646 29428
rect 16716 29316 16772 29372
rect 12562 29260 12572 29316
rect 12628 29260 16660 29316
rect 16716 29260 27916 29316
rect 27972 29260 28364 29316
rect 28420 29260 28430 29316
rect 16604 29204 16660 29260
rect 1922 29148 1932 29204
rect 1988 29148 1998 29204
rect 4946 29148 4956 29204
rect 5012 29148 15148 29204
rect 16604 29148 18396 29204
rect 18452 29148 19180 29204
rect 19236 29148 23548 29204
rect 23604 29148 24332 29204
rect 24388 29148 24398 29204
rect 43362 29148 43372 29204
rect 43428 29148 45276 29204
rect 45332 29148 45342 29204
rect 0 28980 800 29008
rect 1932 28980 1988 29148
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 15092 28980 15148 29148
rect 18946 29036 18956 29092
rect 19012 29036 22540 29092
rect 22596 29036 24668 29092
rect 24724 29036 24734 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 1988 28980
rect 15092 28924 19068 28980
rect 19124 28924 19134 28980
rect 0 28896 800 28924
rect 23202 28700 23212 28756
rect 23268 28700 23772 28756
rect 23828 28700 25900 28756
rect 25956 28700 25966 28756
rect 12898 28588 12908 28644
rect 12964 28588 13916 28644
rect 13972 28588 13982 28644
rect 24994 28588 25004 28644
rect 25060 28588 25564 28644
rect 25620 28588 26572 28644
rect 26628 28588 26638 28644
rect 27906 28588 27916 28644
rect 27972 28588 29148 28644
rect 29204 28588 29214 28644
rect 29474 28588 29484 28644
rect 29540 28588 30268 28644
rect 30324 28588 30334 28644
rect 34402 28588 34412 28644
rect 34468 28588 36988 28644
rect 37044 28588 37054 28644
rect 18498 28476 18508 28532
rect 18564 28476 19068 28532
rect 19124 28476 19134 28532
rect 27682 28476 27692 28532
rect 27748 28476 28140 28532
rect 28196 28476 29372 28532
rect 29428 28476 32732 28532
rect 32788 28476 32798 28532
rect 41010 28476 41020 28532
rect 41076 28476 41580 28532
rect 41636 28476 44492 28532
rect 44548 28476 44558 28532
rect 1698 28364 1708 28420
rect 1764 28364 1774 28420
rect 15092 28364 25676 28420
rect 25732 28364 26124 28420
rect 26180 28364 26908 28420
rect 42018 28364 42028 28420
rect 42084 28364 42812 28420
rect 42868 28364 45164 28420
rect 45220 28364 45230 28420
rect 0 28308 800 28336
rect 1708 28308 1764 28364
rect 0 28252 1764 28308
rect 0 28224 800 28252
rect 15092 28084 15148 28364
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 26852 28084 26908 28364
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 2034 28028 2044 28084
rect 2100 28028 15148 28084
rect 16034 28028 16044 28084
rect 16100 28028 19628 28084
rect 19684 28028 19694 28084
rect 24658 28028 24668 28084
rect 24724 28028 26012 28084
rect 26068 28028 26078 28084
rect 26674 28028 26684 28084
rect 26740 28028 27132 28084
rect 27188 28028 27198 28084
rect 17938 27916 17948 27972
rect 18004 27916 19404 27972
rect 19460 27916 19470 27972
rect 6066 27804 6076 27860
rect 6132 27804 8428 27860
rect 18834 27804 18844 27860
rect 18900 27804 33404 27860
rect 33460 27804 33470 27860
rect 34962 27804 34972 27860
rect 35028 27804 37996 27860
rect 38052 27804 41356 27860
rect 41412 27804 41422 27860
rect 49634 27804 49644 27860
rect 49700 27804 51100 27860
rect 51156 27804 51166 27860
rect 51986 27804 51996 27860
rect 52052 27804 52892 27860
rect 52948 27804 52958 27860
rect 8372 27748 8428 27804
rect 34972 27748 35028 27804
rect 8372 27692 15148 27748
rect 21746 27692 21756 27748
rect 21812 27692 24220 27748
rect 24276 27692 25228 27748
rect 25284 27692 25294 27748
rect 33170 27692 33180 27748
rect 33236 27692 33516 27748
rect 33572 27692 35028 27748
rect 47954 27692 47964 27748
rect 48020 27692 49532 27748
rect 49588 27692 49868 27748
rect 49924 27692 50428 27748
rect 50484 27692 50494 27748
rect 0 27636 800 27664
rect 15092 27636 15148 27692
rect 59200 27636 60000 27664
rect 0 27580 1708 27636
rect 1764 27580 2492 27636
rect 2548 27580 2558 27636
rect 4284 27580 8428 27636
rect 15092 27580 18732 27636
rect 18788 27580 18798 27636
rect 42242 27580 42252 27636
rect 42308 27580 43260 27636
rect 43316 27580 45052 27636
rect 45108 27580 45118 27636
rect 50306 27580 50316 27636
rect 50372 27580 51660 27636
rect 51716 27580 51726 27636
rect 57922 27580 57932 27636
rect 57988 27580 60000 27636
rect 0 27552 800 27580
rect 4284 27524 4340 27580
rect 2034 27468 2044 27524
rect 2100 27468 4340 27524
rect 8372 27524 8428 27580
rect 59200 27552 60000 27580
rect 8372 27468 26908 27524
rect 26964 27468 26974 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 9202 27356 9212 27412
rect 9268 27356 9660 27412
rect 9716 27356 16044 27412
rect 16100 27356 16110 27412
rect 46386 27356 46396 27412
rect 46452 27356 46844 27412
rect 46900 27356 46910 27412
rect 47394 27356 47404 27412
rect 47460 27356 49420 27412
rect 49476 27356 49980 27412
rect 50036 27356 50876 27412
rect 50932 27356 50942 27412
rect 21074 27244 21084 27300
rect 21140 27244 37772 27300
rect 37828 27244 37838 27300
rect 49074 27244 49084 27300
rect 49140 27244 49644 27300
rect 49700 27244 49710 27300
rect 8866 27132 8876 27188
rect 8932 27132 10332 27188
rect 10388 27132 10398 27188
rect 15026 27132 15036 27188
rect 15092 27132 18732 27188
rect 18788 27132 18798 27188
rect 40226 27132 40236 27188
rect 40292 27132 41020 27188
rect 41076 27132 41086 27188
rect 43558 27132 43596 27188
rect 43652 27132 43662 27188
rect 18386 27020 18396 27076
rect 18452 27020 22764 27076
rect 22820 27020 22830 27076
rect 37202 27020 37212 27076
rect 37268 27020 41468 27076
rect 41524 27020 41534 27076
rect 51762 27020 51772 27076
rect 51828 27020 51996 27076
rect 52052 27020 52062 27076
rect 54226 27020 54236 27076
rect 54292 27020 55580 27076
rect 55636 27020 55646 27076
rect 0 26964 800 26992
rect 0 26908 1708 26964
rect 1764 26908 2492 26964
rect 2548 26908 2558 26964
rect 12450 26908 12460 26964
rect 12516 26908 16268 26964
rect 16324 26908 16334 26964
rect 43586 26908 43596 26964
rect 43652 26908 45612 26964
rect 45668 26908 45678 26964
rect 45826 26908 45836 26964
rect 45892 26908 46508 26964
rect 46564 26908 48748 26964
rect 48804 26908 48814 26964
rect 50866 26908 50876 26964
rect 50932 26908 52556 26964
rect 52612 26908 52622 26964
rect 0 26880 800 26908
rect 6290 26796 6300 26852
rect 6356 26796 11396 26852
rect 22866 26796 22876 26852
rect 22932 26796 23548 26852
rect 23604 26796 24332 26852
rect 24388 26796 24398 26852
rect 11340 26740 11396 26796
rect 3332 26684 9436 26740
rect 9492 26684 9502 26740
rect 11330 26684 11340 26740
rect 11396 26684 13468 26740
rect 13524 26684 13534 26740
rect 3332 26516 3388 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 5058 26572 5068 26628
rect 5124 26572 5740 26628
rect 5796 26572 14924 26628
rect 14980 26572 14990 26628
rect 21634 26572 21644 26628
rect 21700 26572 23436 26628
rect 23492 26572 24780 26628
rect 24836 26572 24846 26628
rect 39666 26572 39676 26628
rect 39732 26572 39742 26628
rect 39676 26516 39732 26572
rect 2706 26460 2716 26516
rect 2772 26460 3388 26516
rect 10434 26460 10444 26516
rect 10500 26460 14028 26516
rect 14084 26460 16380 26516
rect 16436 26460 16446 26516
rect 38770 26460 38780 26516
rect 38836 26460 39732 26516
rect 9986 26348 9996 26404
rect 10052 26348 21196 26404
rect 21252 26348 21262 26404
rect 30930 26348 30940 26404
rect 30996 26348 31724 26404
rect 31780 26348 38220 26404
rect 38276 26348 39676 26404
rect 39732 26348 39742 26404
rect 49746 26348 49756 26404
rect 49812 26348 50316 26404
rect 50372 26348 50382 26404
rect 0 26292 800 26320
rect 59200 26292 60000 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 2258 26236 2268 26292
rect 2324 26236 4396 26292
rect 4452 26236 4844 26292
rect 4900 26236 21756 26292
rect 21812 26236 21822 26292
rect 24210 26236 24220 26292
rect 24276 26236 30828 26292
rect 30884 26236 30894 26292
rect 43138 26236 43148 26292
rect 43204 26236 43596 26292
rect 43652 26236 43708 26292
rect 43764 26236 43774 26292
rect 50082 26236 50092 26292
rect 50148 26236 50988 26292
rect 51044 26236 51054 26292
rect 51426 26236 51436 26292
rect 51492 26236 52332 26292
rect 52388 26236 52398 26292
rect 52882 26236 52892 26292
rect 52948 26236 53676 26292
rect 53732 26236 53742 26292
rect 57922 26236 57932 26292
rect 57988 26236 60000 26292
rect 0 26208 800 26236
rect 59200 26208 60000 26236
rect 2370 26124 2380 26180
rect 2436 26124 3164 26180
rect 3220 26124 3230 26180
rect 8194 26124 8204 26180
rect 8260 26124 10780 26180
rect 10836 26124 11340 26180
rect 11396 26124 11406 26180
rect 22866 26124 22876 26180
rect 22932 26124 23996 26180
rect 24052 26124 24062 26180
rect 25890 26124 25900 26180
rect 25956 26124 26684 26180
rect 26740 26124 27468 26180
rect 27524 26124 27534 26180
rect 28998 26124 29036 26180
rect 29092 26124 29102 26180
rect 46498 26124 46508 26180
rect 46564 26124 46956 26180
rect 47012 26124 47022 26180
rect 4274 26012 4284 26068
rect 4340 26012 14476 26068
rect 14532 26012 15036 26068
rect 15092 26012 15102 26068
rect 22082 26012 22092 26068
rect 22148 26012 23436 26068
rect 23492 26012 25340 26068
rect 25396 26012 25406 26068
rect 26114 26012 26124 26068
rect 26180 26012 26908 26068
rect 26964 26012 27244 26068
rect 27300 26012 27310 26068
rect 28354 26012 28364 26068
rect 28420 26012 34188 26068
rect 34244 26012 34254 26068
rect 38658 26012 38668 26068
rect 38724 26012 39228 26068
rect 39284 26012 39294 26068
rect 26124 25956 26180 26012
rect 20626 25900 20636 25956
rect 20692 25900 21420 25956
rect 21476 25900 26180 25956
rect 50530 25900 50540 25956
rect 50596 25900 50876 25956
rect 50932 25900 50942 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 22978 25788 22988 25844
rect 23044 25788 23772 25844
rect 23828 25788 34132 25844
rect 34076 25732 34132 25788
rect 5506 25676 5516 25732
rect 5572 25676 8764 25732
rect 8820 25676 12348 25732
rect 12404 25676 12414 25732
rect 16258 25676 16268 25732
rect 16324 25676 22540 25732
rect 22596 25676 22606 25732
rect 23874 25676 23884 25732
rect 23940 25676 27916 25732
rect 27972 25676 27982 25732
rect 29026 25676 29036 25732
rect 29092 25676 29708 25732
rect 29764 25676 29774 25732
rect 30370 25676 30380 25732
rect 30436 25676 33852 25732
rect 33908 25676 33918 25732
rect 34076 25676 34636 25732
rect 34692 25676 35532 25732
rect 35588 25676 35598 25732
rect 0 25620 800 25648
rect 0 25564 2380 25620
rect 2436 25564 2446 25620
rect 6514 25564 6524 25620
rect 6580 25564 19628 25620
rect 19684 25564 19694 25620
rect 20290 25564 20300 25620
rect 20356 25564 22764 25620
rect 22820 25564 22830 25620
rect 23090 25564 23100 25620
rect 23156 25564 24668 25620
rect 24724 25564 24734 25620
rect 29260 25564 32900 25620
rect 34066 25564 34076 25620
rect 34132 25564 42364 25620
rect 42420 25564 42430 25620
rect 47170 25564 47180 25620
rect 47236 25564 49084 25620
rect 49140 25564 49150 25620
rect 51650 25564 51660 25620
rect 51716 25564 52668 25620
rect 52724 25564 52734 25620
rect 0 25536 800 25564
rect 20300 25508 20356 25564
rect 15092 25452 17836 25508
rect 17892 25452 17902 25508
rect 18162 25452 18172 25508
rect 18228 25452 18732 25508
rect 18788 25452 20356 25508
rect 24770 25452 24780 25508
rect 24836 25452 28252 25508
rect 28308 25452 28318 25508
rect 4386 25340 4396 25396
rect 4452 25340 5180 25396
rect 5236 25340 5246 25396
rect 4162 25228 4172 25284
rect 4228 25228 4732 25284
rect 4788 25228 6300 25284
rect 6356 25228 6366 25284
rect 15092 25172 15148 25452
rect 29260 25396 29316 25564
rect 32844 25508 32900 25564
rect 29474 25452 29484 25508
rect 29540 25452 29550 25508
rect 30706 25452 30716 25508
rect 30772 25452 31500 25508
rect 31556 25452 31566 25508
rect 32834 25452 32844 25508
rect 32900 25452 32910 25508
rect 38994 25452 39004 25508
rect 39060 25452 39070 25508
rect 45154 25452 45164 25508
rect 45220 25452 46284 25508
rect 46340 25452 46844 25508
rect 46900 25452 46910 25508
rect 48850 25452 48860 25508
rect 48916 25452 50204 25508
rect 50260 25452 50652 25508
rect 50708 25452 50718 25508
rect 15362 25340 15372 25396
rect 15428 25340 16044 25396
rect 16100 25340 16110 25396
rect 25778 25340 25788 25396
rect 25844 25340 29316 25396
rect 29484 25284 29540 25452
rect 39004 25284 39060 25452
rect 42354 25340 42364 25396
rect 42420 25340 43372 25396
rect 43428 25340 43438 25396
rect 16594 25228 16604 25284
rect 16660 25228 18564 25284
rect 27682 25228 27692 25284
rect 27748 25228 28700 25284
rect 28756 25228 29540 25284
rect 32050 25228 32060 25284
rect 32116 25228 33740 25284
rect 33796 25228 33806 25284
rect 37314 25228 37324 25284
rect 37380 25228 39060 25284
rect 41234 25228 41244 25284
rect 41300 25228 46508 25284
rect 46564 25228 46574 25284
rect 46946 25228 46956 25284
rect 47012 25228 50764 25284
rect 50820 25228 50830 25284
rect 5954 25116 5964 25172
rect 6020 25116 15148 25172
rect 0 24948 800 24976
rect 18508 24948 18564 25228
rect 20178 25116 20188 25172
rect 20244 25116 23884 25172
rect 23940 25116 23950 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 23314 25004 23324 25060
rect 23380 25004 31948 25060
rect 32004 25004 32014 25060
rect 59200 24948 60000 24976
rect 0 24892 1708 24948
rect 1764 24892 2940 24948
rect 2996 24892 3006 24948
rect 15474 24892 15484 24948
rect 15540 24892 17836 24948
rect 17892 24892 18284 24948
rect 18340 24892 18350 24948
rect 18508 24892 18732 24948
rect 18788 24892 20860 24948
rect 20916 24892 20926 24948
rect 57922 24892 57932 24948
rect 57988 24892 60000 24948
rect 0 24864 800 24892
rect 59200 24864 60000 24892
rect 19170 24780 19180 24836
rect 19236 24780 20972 24836
rect 21028 24780 21038 24836
rect 33618 24780 33628 24836
rect 33684 24780 35196 24836
rect 35252 24780 35262 24836
rect 42578 24780 42588 24836
rect 42644 24780 43372 24836
rect 43428 24780 43438 24836
rect 4274 24668 4284 24724
rect 4340 24668 14140 24724
rect 14196 24668 14924 24724
rect 14980 24668 17388 24724
rect 17444 24668 17454 24724
rect 24994 24668 25004 24724
rect 25060 24668 26012 24724
rect 26068 24668 26078 24724
rect 28018 24668 28028 24724
rect 28084 24668 30828 24724
rect 30884 24668 30894 24724
rect 31266 24668 31276 24724
rect 31332 24668 32060 24724
rect 32116 24668 32126 24724
rect 33282 24668 33292 24724
rect 33348 24668 34300 24724
rect 34356 24668 34366 24724
rect 43474 24668 43484 24724
rect 43540 24668 44716 24724
rect 44772 24668 44782 24724
rect 46274 24668 46284 24724
rect 46340 24668 47068 24724
rect 47124 24668 47134 24724
rect 47954 24668 47964 24724
rect 48020 24668 48972 24724
rect 49028 24668 49038 24724
rect 12226 24556 12236 24612
rect 12292 24556 13916 24612
rect 13972 24556 15260 24612
rect 15316 24556 19068 24612
rect 19124 24556 19134 24612
rect 20402 24556 20412 24612
rect 20468 24556 32620 24612
rect 32676 24556 35644 24612
rect 35700 24556 36428 24612
rect 36484 24556 37100 24612
rect 37156 24556 37166 24612
rect 44370 24556 44380 24612
rect 44436 24556 49308 24612
rect 49364 24556 49374 24612
rect 34860 24500 34916 24556
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 7970 24444 7980 24500
rect 8036 24444 8764 24500
rect 8820 24444 8830 24500
rect 22866 24444 22876 24500
rect 22932 24444 23324 24500
rect 23380 24444 23390 24500
rect 23538 24444 23548 24500
rect 23604 24444 24556 24500
rect 24612 24444 24622 24500
rect 34850 24444 34860 24500
rect 34916 24444 34926 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 17602 24332 17612 24388
rect 17668 24332 18060 24388
rect 18116 24332 25340 24388
rect 25396 24332 25406 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 59200 24276 60000 24304
rect 0 24220 1988 24276
rect 10658 24220 10668 24276
rect 10724 24220 23380 24276
rect 25218 24220 25228 24276
rect 25284 24220 28140 24276
rect 28196 24220 28206 24276
rect 55346 24220 55356 24276
rect 55412 24220 60000 24276
rect 0 24192 800 24220
rect 23324 24164 23380 24220
rect 59200 24192 60000 24220
rect 18274 24108 18284 24164
rect 18340 24108 22876 24164
rect 22932 24108 22942 24164
rect 23314 24108 23324 24164
rect 23380 24108 23390 24164
rect 30034 24108 30044 24164
rect 30100 24108 30716 24164
rect 30772 24108 30782 24164
rect 36194 24108 36204 24164
rect 36260 24108 36988 24164
rect 37044 24108 37054 24164
rect 38612 24108 43148 24164
rect 43204 24108 43214 24164
rect 46834 24108 46844 24164
rect 46900 24108 50428 24164
rect 38612 24052 38668 24108
rect 14364 23996 19292 24052
rect 19348 23996 19358 24052
rect 21410 23996 21420 24052
rect 21476 23996 32788 24052
rect 32946 23996 32956 24052
rect 33012 23996 38668 24052
rect 14364 23940 14420 23996
rect 32732 23940 32788 23996
rect 50372 23940 50428 24108
rect 4274 23884 4284 23940
rect 4340 23884 10108 23940
rect 10164 23884 11228 23940
rect 11284 23884 12572 23940
rect 12628 23884 12638 23940
rect 14354 23884 14364 23940
rect 14420 23884 14430 23940
rect 14578 23884 14588 23940
rect 14644 23884 16492 23940
rect 16548 23884 16558 23940
rect 18610 23884 18620 23940
rect 18676 23884 19852 23940
rect 19908 23884 19918 23940
rect 22978 23884 22988 23940
rect 23044 23884 27132 23940
rect 27188 23884 27198 23940
rect 30258 23884 30268 23940
rect 30324 23884 31164 23940
rect 31220 23884 31230 23940
rect 32732 23884 35756 23940
rect 35812 23884 36204 23940
rect 36260 23884 36270 23940
rect 36754 23884 36764 23940
rect 36820 23884 38780 23940
rect 38836 23884 38846 23940
rect 47170 23884 47180 23940
rect 47236 23884 48188 23940
rect 48244 23884 48748 23940
rect 48804 23884 48814 23940
rect 50372 23884 55580 23940
rect 55636 23884 55646 23940
rect 36204 23828 36260 23884
rect 16146 23772 16156 23828
rect 16212 23772 22204 23828
rect 22260 23772 22270 23828
rect 22866 23772 22876 23828
rect 22932 23772 23772 23828
rect 23828 23772 23838 23828
rect 24994 23772 25004 23828
rect 25060 23772 25564 23828
rect 25620 23772 26460 23828
rect 26516 23772 26684 23828
rect 26740 23772 26750 23828
rect 27570 23772 27580 23828
rect 27636 23772 33292 23828
rect 33348 23772 33964 23828
rect 34020 23772 34030 23828
rect 34738 23772 34748 23828
rect 34804 23772 35252 23828
rect 35308 23772 35318 23828
rect 36204 23772 40348 23828
rect 40404 23772 40414 23828
rect 7298 23660 7308 23716
rect 7364 23660 9100 23716
rect 9156 23660 9166 23716
rect 20962 23660 20972 23716
rect 21028 23660 23100 23716
rect 23156 23660 23166 23716
rect 24882 23660 24892 23716
rect 24948 23660 25340 23716
rect 25396 23660 25406 23716
rect 29474 23660 29484 23716
rect 29540 23660 30268 23716
rect 30324 23660 30334 23716
rect 30594 23660 30604 23716
rect 30660 23660 37828 23716
rect 42018 23660 42028 23716
rect 42084 23660 42700 23716
rect 42756 23660 42766 23716
rect 0 23604 800 23632
rect 37772 23604 37828 23660
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 16482 23548 16492 23604
rect 16548 23548 18620 23604
rect 18676 23548 18686 23604
rect 21942 23548 21980 23604
rect 22036 23548 22046 23604
rect 22194 23548 22204 23604
rect 22260 23548 31724 23604
rect 31780 23548 31790 23604
rect 34178 23548 34188 23604
rect 34244 23548 35644 23604
rect 35700 23548 35710 23604
rect 36866 23548 36876 23604
rect 36932 23548 37100 23604
rect 37156 23548 37166 23604
rect 37762 23548 37772 23604
rect 37828 23548 37838 23604
rect 38546 23548 38556 23604
rect 38612 23548 47964 23604
rect 48020 23548 48030 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 11666 23436 11676 23492
rect 11732 23436 13860 23492
rect 14914 23436 14924 23492
rect 14980 23436 16268 23492
rect 16324 23436 16334 23492
rect 28354 23436 28364 23492
rect 28420 23436 34972 23492
rect 35028 23436 35038 23492
rect 35410 23436 35420 23492
rect 35476 23436 36204 23492
rect 36260 23436 36270 23492
rect 44258 23436 44268 23492
rect 44324 23436 44940 23492
rect 44996 23436 45006 23492
rect 51426 23436 51436 23492
rect 51492 23436 52780 23492
rect 52836 23436 52846 23492
rect 13804 23380 13860 23436
rect 4162 23324 4172 23380
rect 4228 23324 8764 23380
rect 8820 23324 9548 23380
rect 9604 23324 9614 23380
rect 11890 23324 11900 23380
rect 11956 23324 12796 23380
rect 12852 23324 13580 23380
rect 13636 23324 13646 23380
rect 13804 23324 24556 23380
rect 24612 23324 24622 23380
rect 25666 23324 25676 23380
rect 25732 23324 26124 23380
rect 26180 23324 26908 23380
rect 26964 23324 28140 23380
rect 28196 23324 28206 23380
rect 34402 23324 34412 23380
rect 34468 23324 45388 23380
rect 45444 23324 45454 23380
rect 50194 23324 50204 23380
rect 50260 23324 51100 23380
rect 51156 23324 51884 23380
rect 51940 23324 51950 23380
rect 52210 23324 52220 23380
rect 52276 23324 52892 23380
rect 52948 23324 52958 23380
rect 4274 23212 4284 23268
rect 4340 23212 7868 23268
rect 7924 23212 8876 23268
rect 8932 23212 8942 23268
rect 12002 23212 12012 23268
rect 12068 23212 12684 23268
rect 12740 23212 16716 23268
rect 16772 23212 26908 23268
rect 27458 23212 27468 23268
rect 27524 23212 28476 23268
rect 28532 23212 28542 23268
rect 31826 23212 31836 23268
rect 31892 23212 32508 23268
rect 32564 23212 32574 23268
rect 35858 23212 35868 23268
rect 35924 23212 37996 23268
rect 38052 23212 38062 23268
rect 40002 23212 40012 23268
rect 40068 23212 41020 23268
rect 41076 23212 41086 23268
rect 41794 23212 41804 23268
rect 41860 23212 42812 23268
rect 42868 23212 43148 23268
rect 43204 23212 43214 23268
rect 47618 23212 47628 23268
rect 47684 23212 51212 23268
rect 51268 23212 51660 23268
rect 51716 23212 51726 23268
rect 8306 23100 8316 23156
rect 8372 23100 9324 23156
rect 9380 23100 10556 23156
rect 10612 23100 10622 23156
rect 13906 23100 13916 23156
rect 13972 23100 16268 23156
rect 16324 23100 16334 23156
rect 20290 23100 20300 23156
rect 20356 23100 21420 23156
rect 21476 23100 21486 23156
rect 12898 22988 12908 23044
rect 12964 22988 22540 23044
rect 22596 22988 22606 23044
rect 26086 22988 26124 23044
rect 26180 22988 26684 23044
rect 26740 22988 26750 23044
rect 0 22932 800 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 24322 22876 24332 22932
rect 24388 22876 25340 22932
rect 25396 22876 25406 22932
rect 0 22848 800 22876
rect 26852 22820 26908 23212
rect 27010 23100 27020 23156
rect 27076 23100 27692 23156
rect 27748 23100 28364 23156
rect 28420 23100 28430 23156
rect 31490 23100 31500 23156
rect 31556 23100 34300 23156
rect 34356 23100 34366 23156
rect 40114 23100 40124 23156
rect 40180 23100 40908 23156
rect 40964 23100 40974 23156
rect 43586 23100 43596 23156
rect 43652 23100 44156 23156
rect 44212 23100 44222 23156
rect 30370 22988 30380 23044
rect 30436 22988 32172 23044
rect 32228 22988 32238 23044
rect 33730 22988 33740 23044
rect 33796 22988 34524 23044
rect 34580 22988 34590 23044
rect 35186 22988 35196 23044
rect 35252 22988 38332 23044
rect 38388 22988 39004 23044
rect 39060 22988 39070 23044
rect 42130 22988 42140 23044
rect 42196 22988 47292 23044
rect 47348 22988 47358 23044
rect 28018 22876 28028 22932
rect 28084 22876 30268 22932
rect 30324 22876 30334 22932
rect 31042 22876 31052 22932
rect 31108 22876 39116 22932
rect 39172 22876 39676 22932
rect 39732 22876 39742 22932
rect 26852 22764 28364 22820
rect 28420 22764 28430 22820
rect 37538 22764 37548 22820
rect 37604 22764 38220 22820
rect 38276 22764 38286 22820
rect 39218 22764 39228 22820
rect 39284 22764 40124 22820
rect 40180 22764 41020 22820
rect 41076 22764 41916 22820
rect 41972 22764 42364 22820
rect 42420 22764 42430 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19506 22652 19516 22708
rect 19572 22652 20076 22708
rect 20132 22652 26908 22708
rect 28242 22652 28252 22708
rect 28308 22652 31388 22708
rect 31444 22652 32508 22708
rect 32564 22652 32574 22708
rect 36194 22652 36204 22708
rect 36260 22652 39004 22708
rect 39060 22652 39788 22708
rect 39844 22652 40796 22708
rect 40852 22652 40862 22708
rect 47964 22652 52892 22708
rect 52948 22652 52958 22708
rect 26852 22596 26908 22652
rect 47964 22596 48020 22652
rect 26852 22540 31108 22596
rect 31266 22540 31276 22596
rect 31332 22540 44492 22596
rect 44548 22540 45388 22596
rect 45444 22540 45454 22596
rect 47954 22540 47964 22596
rect 48020 22540 48030 22596
rect 31052 22484 31108 22540
rect 1922 22428 1932 22484
rect 1988 22428 1998 22484
rect 10882 22428 10892 22484
rect 10948 22428 13020 22484
rect 13076 22428 13086 22484
rect 15362 22428 15372 22484
rect 15428 22428 17164 22484
rect 17220 22428 17230 22484
rect 20524 22428 21980 22484
rect 22036 22428 22046 22484
rect 26898 22428 26908 22484
rect 26964 22428 27804 22484
rect 27860 22428 27870 22484
rect 31052 22428 33628 22484
rect 33684 22428 35084 22484
rect 35140 22428 35150 22484
rect 38098 22428 38108 22484
rect 38164 22428 43708 22484
rect 43764 22428 43774 22484
rect 47282 22428 47292 22484
rect 47348 22428 47740 22484
rect 47796 22428 47806 22484
rect 50372 22428 50876 22484
rect 50932 22428 50942 22484
rect 0 22260 800 22288
rect 1932 22260 1988 22428
rect 20524 22372 20580 22428
rect 50372 22372 50428 22428
rect 8978 22316 8988 22372
rect 9044 22316 9660 22372
rect 9716 22316 11564 22372
rect 11620 22316 11630 22372
rect 13906 22316 13916 22372
rect 13972 22316 14588 22372
rect 14644 22316 14654 22372
rect 16370 22316 16380 22372
rect 16436 22316 17276 22372
rect 17332 22316 17342 22372
rect 19058 22316 19068 22372
rect 19124 22316 20524 22372
rect 20580 22316 20590 22372
rect 20850 22316 20860 22372
rect 20916 22316 21532 22372
rect 21588 22316 24780 22372
rect 24836 22316 24846 22372
rect 26562 22316 26572 22372
rect 26628 22316 28252 22372
rect 28308 22316 29932 22372
rect 29988 22316 29998 22372
rect 43810 22316 43820 22372
rect 43876 22316 50204 22372
rect 50260 22316 50428 22372
rect 53106 22316 53116 22372
rect 53172 22316 54460 22372
rect 54516 22316 54526 22372
rect 0 22204 1988 22260
rect 6290 22204 6300 22260
rect 6356 22204 9772 22260
rect 9828 22204 9838 22260
rect 15138 22204 15148 22260
rect 15204 22204 15820 22260
rect 15876 22204 18284 22260
rect 18340 22204 19292 22260
rect 19348 22204 19358 22260
rect 24434 22204 24444 22260
rect 24500 22204 25452 22260
rect 25508 22204 27132 22260
rect 27188 22204 27198 22260
rect 29138 22204 29148 22260
rect 29204 22204 30044 22260
rect 30100 22204 30940 22260
rect 30996 22204 31006 22260
rect 53218 22204 53228 22260
rect 53284 22204 54236 22260
rect 54292 22204 54302 22260
rect 0 22176 800 22204
rect 6850 22092 6860 22148
rect 6916 22092 8428 22148
rect 8484 22092 10220 22148
rect 10276 22092 10780 22148
rect 10836 22092 11228 22148
rect 11284 22092 11294 22148
rect 11778 22092 11788 22148
rect 11844 22092 12348 22148
rect 12404 22092 12414 22148
rect 12870 22092 12908 22148
rect 12964 22092 12974 22148
rect 13458 22092 13468 22148
rect 13524 22092 20244 22148
rect 25218 22092 25228 22148
rect 25284 22092 29708 22148
rect 29764 22092 29774 22148
rect 35410 22092 35420 22148
rect 35476 22092 41132 22148
rect 41188 22092 41198 22148
rect 43362 22092 43372 22148
rect 43428 22092 43932 22148
rect 43988 22092 45500 22148
rect 45556 22092 45566 22148
rect 50428 22092 50652 22148
rect 50708 22092 50718 22148
rect 12908 22036 12964 22092
rect 20188 22036 20244 22092
rect 12908 21980 16044 22036
rect 16100 21980 17892 22036
rect 20188 21980 27132 22036
rect 27188 21980 27198 22036
rect 30678 21980 30716 22036
rect 30772 21980 30782 22036
rect 37650 21980 37660 22036
rect 37716 21980 38108 22036
rect 38164 21980 38174 22036
rect 46050 21980 46060 22036
rect 46116 21980 46284 22036
rect 46340 21980 47404 22036
rect 47460 21980 47470 22036
rect 11106 21868 11116 21924
rect 11172 21868 11900 21924
rect 11956 21868 11966 21924
rect 16706 21868 16716 21924
rect 16772 21868 17500 21924
rect 17556 21868 17566 21924
rect 17836 21812 17892 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 21644 21868 22428 21924
rect 22484 21868 22494 21924
rect 24658 21868 24668 21924
rect 24724 21868 25116 21924
rect 25172 21868 25182 21924
rect 27794 21868 27804 21924
rect 27860 21868 39452 21924
rect 39508 21868 39518 21924
rect 42802 21868 42812 21924
rect 42868 21868 43036 21924
rect 43092 21868 43596 21924
rect 43652 21868 44156 21924
rect 44212 21868 44222 21924
rect 44930 21868 44940 21924
rect 44996 21868 45948 21924
rect 46004 21868 46014 21924
rect 21644 21812 21700 21868
rect 50428 21812 50484 22092
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4274 21756 4284 21812
rect 4340 21756 6748 21812
rect 6804 21756 7420 21812
rect 7476 21756 7980 21812
rect 8036 21756 8046 21812
rect 14242 21756 14252 21812
rect 14308 21756 16492 21812
rect 16548 21756 16558 21812
rect 17836 21756 21644 21812
rect 21700 21756 21710 21812
rect 22306 21756 22316 21812
rect 22372 21756 22764 21812
rect 22820 21756 22830 21812
rect 22978 21756 22988 21812
rect 23044 21756 25340 21812
rect 25396 21756 25406 21812
rect 27682 21756 27692 21812
rect 27748 21756 33404 21812
rect 33460 21756 33470 21812
rect 34290 21756 34300 21812
rect 34356 21756 35980 21812
rect 36036 21756 36046 21812
rect 42130 21756 42140 21812
rect 42196 21756 44828 21812
rect 44884 21756 44894 21812
rect 50428 21756 50540 21812
rect 50596 21756 50606 21812
rect 15474 21644 15484 21700
rect 15540 21644 18060 21700
rect 18116 21644 18126 21700
rect 18498 21644 18508 21700
rect 18564 21644 19404 21700
rect 19460 21644 19470 21700
rect 20738 21644 20748 21700
rect 20804 21644 21868 21700
rect 21924 21644 21934 21700
rect 22092 21644 26236 21700
rect 26292 21644 26302 21700
rect 31378 21644 31388 21700
rect 31444 21644 33068 21700
rect 33124 21644 33740 21700
rect 33796 21644 34748 21700
rect 34804 21644 34814 21700
rect 36866 21644 36876 21700
rect 36932 21644 49420 21700
rect 49476 21644 49486 21700
rect 0 21588 800 21616
rect 22092 21588 22148 21644
rect 0 21532 1988 21588
rect 5954 21532 5964 21588
rect 6020 21532 6972 21588
rect 7028 21532 7038 21588
rect 14476 21532 14980 21588
rect 15138 21532 15148 21588
rect 15204 21532 16044 21588
rect 16100 21532 17948 21588
rect 18004 21532 18014 21588
rect 20514 21532 20524 21588
rect 20580 21532 22148 21588
rect 22204 21532 24332 21588
rect 24388 21532 24398 21588
rect 24658 21532 24668 21588
rect 24724 21532 25340 21588
rect 25396 21532 25788 21588
rect 25844 21532 25854 21588
rect 29362 21532 29372 21588
rect 29428 21532 30828 21588
rect 30884 21532 30894 21588
rect 42802 21532 42812 21588
rect 42868 21532 43484 21588
rect 43540 21532 43550 21588
rect 46834 21532 46844 21588
rect 46900 21532 47404 21588
rect 47460 21532 47470 21588
rect 0 21504 800 21532
rect 1932 21476 1988 21532
rect 14476 21476 14532 21532
rect 14924 21476 14980 21532
rect 22204 21476 22260 21532
rect 1922 21420 1932 21476
rect 1988 21420 1998 21476
rect 11330 21420 11340 21476
rect 11396 21420 13244 21476
rect 13300 21420 13310 21476
rect 14466 21420 14476 21476
rect 14532 21420 14542 21476
rect 14690 21420 14700 21476
rect 14756 21420 14766 21476
rect 14924 21420 22260 21476
rect 24210 21420 24220 21476
rect 24276 21420 26124 21476
rect 26180 21420 26190 21476
rect 30258 21420 30268 21476
rect 30324 21420 31052 21476
rect 31108 21420 31118 21476
rect 40450 21420 40460 21476
rect 40516 21420 41244 21476
rect 41300 21420 41468 21476
rect 41524 21420 42252 21476
rect 42308 21420 42318 21476
rect 53554 21420 53564 21476
rect 53620 21420 54460 21476
rect 54516 21420 54526 21476
rect 14700 21364 14756 21420
rect 14700 21308 16268 21364
rect 16324 21308 18620 21364
rect 18676 21308 19628 21364
rect 19684 21308 19694 21364
rect 24518 21308 24556 21364
rect 24612 21308 27580 21364
rect 27636 21308 27646 21364
rect 31266 21308 31276 21364
rect 31332 21308 37212 21364
rect 37268 21308 37278 21364
rect 38434 21308 38444 21364
rect 38500 21308 38668 21364
rect 41906 21308 41916 21364
rect 41972 21308 42476 21364
rect 42532 21308 42542 21364
rect 46162 21308 46172 21364
rect 46228 21308 51548 21364
rect 51604 21308 51614 21364
rect 17378 21196 17388 21252
rect 17444 21196 22652 21252
rect 22708 21196 23100 21252
rect 23156 21196 23166 21252
rect 23762 21196 23772 21252
rect 23828 21196 25116 21252
rect 25172 21196 25182 21252
rect 25890 21196 25900 21252
rect 25956 21196 29372 21252
rect 29428 21196 29438 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 38612 21140 38668 21308
rect 23874 21084 23884 21140
rect 23940 21084 27916 21140
rect 27972 21084 28308 21140
rect 31714 21084 31724 21140
rect 31780 21084 32284 21140
rect 32340 21084 32350 21140
rect 38612 21084 49196 21140
rect 49252 21084 49262 21140
rect 18722 20972 18732 21028
rect 18788 20972 20524 21028
rect 20580 20972 20590 21028
rect 22418 20972 22428 21028
rect 22484 20972 22876 21028
rect 22932 20972 23548 21028
rect 23604 20972 28028 21028
rect 28084 20972 28094 21028
rect 28252 20916 28308 21084
rect 30146 20972 30156 21028
rect 30212 20972 30828 21028
rect 30884 20972 34188 21028
rect 34244 20972 34254 21028
rect 59200 20916 60000 20944
rect 12450 20860 12460 20916
rect 12516 20860 13468 20916
rect 13524 20860 13534 20916
rect 13682 20860 13692 20916
rect 13748 20860 13804 20916
rect 13860 20860 23772 20916
rect 23828 20860 24108 20916
rect 24164 20860 24174 20916
rect 24332 20860 27244 20916
rect 27300 20860 27310 20916
rect 28252 20860 29596 20916
rect 29652 20860 32844 20916
rect 32900 20860 32910 20916
rect 36978 20860 36988 20916
rect 37044 20860 38220 20916
rect 38276 20860 38286 20916
rect 50530 20860 50540 20916
rect 50596 20860 51212 20916
rect 51268 20860 51278 20916
rect 51762 20860 51772 20916
rect 51828 20860 53340 20916
rect 53396 20860 53406 20916
rect 57922 20860 57932 20916
rect 57988 20860 60000 20916
rect 24332 20804 24388 20860
rect 59200 20832 60000 20860
rect 5842 20748 5852 20804
rect 5908 20748 7868 20804
rect 7924 20748 7934 20804
rect 17164 20748 20524 20804
rect 20580 20748 20590 20804
rect 22418 20748 22428 20804
rect 22484 20748 24388 20804
rect 26562 20748 26572 20804
rect 26628 20748 33628 20804
rect 33684 20748 33694 20804
rect 35858 20748 35868 20804
rect 35924 20748 37996 20804
rect 38052 20748 38062 20804
rect 17164 20692 17220 20748
rect 10994 20636 11004 20692
rect 11060 20636 11564 20692
rect 11620 20636 17164 20692
rect 17220 20636 17230 20692
rect 19730 20636 19740 20692
rect 19796 20636 21532 20692
rect 21588 20636 21598 20692
rect 25666 20636 25676 20692
rect 25732 20636 31164 20692
rect 31220 20636 31230 20692
rect 34066 20636 34076 20692
rect 34132 20636 35084 20692
rect 35140 20636 35150 20692
rect 36082 20636 36092 20692
rect 36148 20636 40572 20692
rect 40628 20636 41580 20692
rect 41636 20636 42140 20692
rect 42196 20636 42206 20692
rect 46386 20636 46396 20692
rect 46452 20636 47740 20692
rect 47796 20636 47806 20692
rect 8866 20524 8876 20580
rect 8932 20524 9772 20580
rect 9828 20524 10668 20580
rect 10724 20524 10734 20580
rect 17826 20524 17836 20580
rect 17892 20524 18620 20580
rect 18676 20524 18686 20580
rect 19170 20524 19180 20580
rect 19236 20524 24892 20580
rect 24948 20524 24958 20580
rect 26226 20524 26236 20580
rect 26292 20524 26572 20580
rect 26628 20524 27356 20580
rect 27412 20524 27422 20580
rect 28018 20524 28028 20580
rect 28084 20524 28364 20580
rect 28420 20524 28430 20580
rect 29922 20524 29932 20580
rect 29988 20524 30380 20580
rect 30436 20524 31388 20580
rect 31444 20524 31454 20580
rect 45378 20524 45388 20580
rect 45444 20524 46172 20580
rect 46228 20524 46238 20580
rect 49410 20524 49420 20580
rect 49476 20524 50540 20580
rect 50596 20524 50606 20580
rect 3266 20412 3276 20468
rect 3332 20412 13580 20468
rect 13636 20412 18508 20468
rect 18564 20412 19628 20468
rect 19684 20412 19694 20468
rect 21410 20412 21420 20468
rect 21476 20412 22316 20468
rect 22372 20412 23324 20468
rect 23380 20412 23390 20468
rect 27906 20412 27916 20468
rect 27972 20412 28812 20468
rect 28868 20412 28878 20468
rect 29362 20412 29372 20468
rect 29428 20412 31836 20468
rect 31892 20412 31902 20468
rect 41682 20412 41692 20468
rect 41748 20412 42812 20468
rect 42868 20412 42878 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 6290 20300 6300 20356
rect 6356 20300 14028 20356
rect 14084 20300 14094 20356
rect 14802 20300 14812 20356
rect 14868 20300 17388 20356
rect 17444 20300 17454 20356
rect 18386 20300 18396 20356
rect 18452 20300 18462 20356
rect 21746 20300 21756 20356
rect 21812 20300 30492 20356
rect 30548 20300 30558 20356
rect 33282 20300 33292 20356
rect 33348 20300 34468 20356
rect 18396 20244 18452 20300
rect 34412 20244 34468 20300
rect 8194 20188 8204 20244
rect 8260 20188 12012 20244
rect 12068 20188 15484 20244
rect 15540 20188 15550 20244
rect 15698 20188 15708 20244
rect 15764 20188 16492 20244
rect 16548 20188 16558 20244
rect 16828 20188 19180 20244
rect 19236 20188 19246 20244
rect 23202 20188 23212 20244
rect 23268 20188 23772 20244
rect 23828 20188 23838 20244
rect 24098 20188 24108 20244
rect 24164 20188 28588 20244
rect 28644 20188 28654 20244
rect 30258 20188 30268 20244
rect 30324 20188 30334 20244
rect 31154 20188 31164 20244
rect 31220 20188 33964 20244
rect 34020 20188 34030 20244
rect 34402 20188 34412 20244
rect 34468 20188 34478 20244
rect 45276 20188 46620 20244
rect 46676 20188 46686 20244
rect 16828 20132 16884 20188
rect 30268 20132 30324 20188
rect 45276 20132 45332 20188
rect 8642 20076 8652 20132
rect 8708 20076 9996 20132
rect 10052 20076 12348 20132
rect 12404 20076 12414 20132
rect 16818 20076 16828 20132
rect 16884 20076 16894 20132
rect 18386 20076 18396 20132
rect 18452 20076 21308 20132
rect 21364 20076 21374 20132
rect 23650 20076 23660 20132
rect 23716 20076 31836 20132
rect 31892 20076 31902 20132
rect 33730 20076 33740 20132
rect 33796 20076 34300 20132
rect 34356 20076 34636 20132
rect 34692 20076 34702 20132
rect 35858 20076 35868 20132
rect 35924 20076 36540 20132
rect 36596 20076 36606 20132
rect 37426 20076 37436 20132
rect 37492 20076 45332 20132
rect 46834 20076 46844 20132
rect 46900 20076 49644 20132
rect 49700 20076 49710 20132
rect 6402 19964 6412 20020
rect 6468 19964 7084 20020
rect 7140 19964 7150 20020
rect 16146 19964 16156 20020
rect 16212 19964 16604 20020
rect 16660 19964 16670 20020
rect 16930 19964 16940 20020
rect 16996 19964 17724 20020
rect 17780 19964 17790 20020
rect 20738 19964 20748 20020
rect 20804 19964 21532 20020
rect 21588 19964 21598 20020
rect 25106 19964 25116 20020
rect 25172 19964 26684 20020
rect 26740 19964 32396 20020
rect 32452 19964 34412 20020
rect 34468 19964 34478 20020
rect 35252 19964 35756 20020
rect 35812 19964 35822 20020
rect 36194 19964 36204 20020
rect 36260 19964 37996 20020
rect 38052 19964 38062 20020
rect 45266 19964 45276 20020
rect 45332 19964 45500 20020
rect 45556 19964 45566 20020
rect 6066 19852 6076 19908
rect 6132 19852 6748 19908
rect 6804 19852 6814 19908
rect 11890 19852 11900 19908
rect 11956 19852 14588 19908
rect 14644 19852 14654 19908
rect 20626 19852 20636 19908
rect 20692 19852 24108 19908
rect 24164 19852 24174 19908
rect 30930 19852 30940 19908
rect 30996 19852 32172 19908
rect 32228 19852 32238 19908
rect 35252 19796 35308 19964
rect 35410 19852 35420 19908
rect 35476 19852 36876 19908
rect 36932 19852 36942 19908
rect 41794 19852 41804 19908
rect 41860 19852 46956 19908
rect 47012 19852 47022 19908
rect 7634 19740 7644 19796
rect 7700 19740 10668 19796
rect 10724 19740 10734 19796
rect 10994 19740 11004 19796
rect 11060 19740 14476 19796
rect 14532 19740 14542 19796
rect 24322 19740 24332 19796
rect 24388 19740 25676 19796
rect 25732 19740 25742 19796
rect 30146 19740 30156 19796
rect 30212 19740 35308 19796
rect 35634 19740 35644 19796
rect 35700 19740 37212 19796
rect 37268 19740 37278 19796
rect 19058 19628 19068 19684
rect 19124 19628 21308 19684
rect 21364 19628 24780 19684
rect 24836 19628 30604 19684
rect 30660 19628 30670 19684
rect 38434 19628 38444 19684
rect 38500 19628 40012 19684
rect 40068 19628 40078 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 22082 19516 22092 19572
rect 22148 19516 22764 19572
rect 22820 19516 25340 19572
rect 25396 19516 25406 19572
rect 27346 19516 27356 19572
rect 27412 19516 28924 19572
rect 28980 19516 28990 19572
rect 15138 19404 15148 19460
rect 15204 19404 15596 19460
rect 15652 19404 18844 19460
rect 18900 19404 19068 19460
rect 19124 19404 19134 19460
rect 23650 19404 23660 19460
rect 23716 19404 24332 19460
rect 24388 19404 24398 19460
rect 26786 19404 26796 19460
rect 26852 19404 28140 19460
rect 28196 19404 28206 19460
rect 30370 19404 30380 19460
rect 30436 19404 30446 19460
rect 32050 19404 32060 19460
rect 32116 19404 35868 19460
rect 35924 19404 36316 19460
rect 36372 19404 36382 19460
rect 26796 19348 26852 19404
rect 21522 19292 21532 19348
rect 21588 19292 22428 19348
rect 22484 19292 25340 19348
rect 25396 19292 26852 19348
rect 30380 19348 30436 19404
rect 30380 19292 43932 19348
rect 43988 19292 43998 19348
rect 10098 19180 10108 19236
rect 10164 19180 20076 19236
rect 20132 19180 26460 19236
rect 26516 19180 26526 19236
rect 26674 19180 26684 19236
rect 26740 19180 29484 19236
rect 29540 19180 29550 19236
rect 31490 19180 31500 19236
rect 31556 19180 32956 19236
rect 33012 19180 34300 19236
rect 34356 19180 34366 19236
rect 46610 19180 46620 19236
rect 46676 19180 47628 19236
rect 47684 19180 47694 19236
rect 51874 19180 51884 19236
rect 51940 19180 53228 19236
rect 53284 19180 53294 19236
rect 7410 19068 7420 19124
rect 7476 19068 7980 19124
rect 8036 19068 8046 19124
rect 16146 19068 16156 19124
rect 16212 19068 19740 19124
rect 19796 19068 20412 19124
rect 20468 19068 20478 19124
rect 25778 19068 25788 19124
rect 25844 19068 27132 19124
rect 27188 19068 27692 19124
rect 27748 19068 27758 19124
rect 1698 18956 1708 19012
rect 1764 18956 1774 19012
rect 8642 18956 8652 19012
rect 8708 18956 9212 19012
rect 9268 18956 9660 19012
rect 9716 18956 11564 19012
rect 11620 18956 12908 19012
rect 12964 18956 20748 19012
rect 20804 18956 21756 19012
rect 21812 18956 24332 19012
rect 24388 18956 24398 19012
rect 28018 18956 28028 19012
rect 28084 18956 30268 19012
rect 30324 18956 30334 19012
rect 36530 18956 36540 19012
rect 36596 18956 37436 19012
rect 37492 18956 38220 19012
rect 38276 18956 38286 19012
rect 42130 18956 42140 19012
rect 42196 18956 46060 19012
rect 46116 18956 46126 19012
rect 46274 18956 46284 19012
rect 46340 18956 46956 19012
rect 47012 18956 47022 19012
rect 50372 18956 50540 19012
rect 50596 18956 52892 19012
rect 52948 18956 52958 19012
rect 0 18900 800 18928
rect 1708 18900 1764 18956
rect 0 18844 1764 18900
rect 9090 18844 9100 18900
rect 9156 18844 11340 18900
rect 11396 18844 18172 18900
rect 18228 18844 18238 18900
rect 23650 18844 23660 18900
rect 23716 18844 25900 18900
rect 25956 18844 25966 18900
rect 37090 18844 37100 18900
rect 37156 18844 37884 18900
rect 37940 18844 37950 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 10770 18732 10780 18788
rect 10836 18732 11340 18788
rect 11396 18732 11406 18788
rect 12898 18732 12908 18788
rect 12964 18732 16436 18788
rect 17490 18732 17500 18788
rect 17556 18732 18732 18788
rect 18788 18732 18798 18788
rect 26338 18732 26348 18788
rect 26404 18732 28140 18788
rect 28196 18732 28206 18788
rect 7858 18620 7868 18676
rect 7924 18620 8204 18676
rect 8260 18620 8270 18676
rect 12338 18620 12348 18676
rect 12404 18620 13692 18676
rect 13748 18620 13758 18676
rect 16380 18564 16436 18732
rect 16706 18620 16716 18676
rect 16772 18620 16940 18676
rect 16996 18620 22036 18676
rect 24434 18620 24444 18676
rect 24500 18620 25788 18676
rect 25844 18620 25854 18676
rect 27682 18620 27692 18676
rect 27748 18620 29036 18676
rect 29092 18620 29102 18676
rect 29586 18620 29596 18676
rect 29652 18620 33180 18676
rect 33236 18620 33246 18676
rect 34514 18620 34524 18676
rect 34580 18620 34860 18676
rect 34916 18620 35756 18676
rect 35812 18620 35822 18676
rect 43586 18620 43596 18676
rect 43652 18620 45724 18676
rect 45780 18620 45790 18676
rect 5730 18508 5740 18564
rect 5796 18508 6748 18564
rect 6804 18508 6814 18564
rect 12786 18508 12796 18564
rect 12852 18508 16156 18564
rect 16212 18508 16222 18564
rect 16370 18508 16380 18564
rect 16436 18508 17948 18564
rect 18004 18508 21308 18564
rect 21364 18508 21374 18564
rect 21980 18452 22036 18620
rect 25890 18508 25900 18564
rect 25956 18508 28364 18564
rect 28420 18508 28924 18564
rect 28980 18508 28990 18564
rect 44818 18508 44828 18564
rect 44884 18508 47068 18564
rect 47124 18508 47134 18564
rect 50372 18452 50428 18956
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 53218 18508 53228 18564
rect 53284 18508 55132 18564
rect 55188 18508 55198 18564
rect 6514 18396 6524 18452
rect 6580 18396 6972 18452
rect 7028 18396 7038 18452
rect 7186 18396 7196 18452
rect 7252 18396 8764 18452
rect 8820 18396 9884 18452
rect 9940 18396 9950 18452
rect 11106 18396 11116 18452
rect 11172 18396 11676 18452
rect 11732 18396 11742 18452
rect 13682 18396 13692 18452
rect 13748 18396 14476 18452
rect 14532 18396 14542 18452
rect 14802 18396 14812 18452
rect 14868 18396 16044 18452
rect 16100 18396 16110 18452
rect 20402 18396 20412 18452
rect 20468 18396 20748 18452
rect 20804 18396 20814 18452
rect 21942 18396 21980 18452
rect 22036 18396 22046 18452
rect 25554 18396 25564 18452
rect 25620 18396 25630 18452
rect 26786 18396 26796 18452
rect 26852 18396 27580 18452
rect 27636 18396 27646 18452
rect 30482 18396 30492 18452
rect 30548 18396 35196 18452
rect 35252 18396 35262 18452
rect 37986 18396 37996 18452
rect 38052 18396 39788 18452
rect 39844 18396 39854 18452
rect 41794 18396 41804 18452
rect 41860 18396 42588 18452
rect 42644 18396 43372 18452
rect 43428 18396 43438 18452
rect 47170 18396 47180 18452
rect 47236 18396 48972 18452
rect 49028 18396 49038 18452
rect 49522 18396 49532 18452
rect 49588 18396 50428 18452
rect 51090 18396 51100 18452
rect 51156 18396 51660 18452
rect 51716 18396 52668 18452
rect 52724 18396 53564 18452
rect 53620 18396 53630 18452
rect 6972 18340 7028 18396
rect 6972 18284 9548 18340
rect 9604 18284 9614 18340
rect 10546 18284 10556 18340
rect 10612 18284 12348 18340
rect 12404 18284 12414 18340
rect 13692 18228 13748 18396
rect 25564 18340 25620 18396
rect 17826 18284 17836 18340
rect 17892 18284 20524 18340
rect 20580 18284 25620 18340
rect 28130 18284 28140 18340
rect 28196 18284 32172 18340
rect 32228 18284 32238 18340
rect 33852 18284 37044 18340
rect 7970 18172 7980 18228
rect 8036 18172 13748 18228
rect 17836 18116 17892 18284
rect 33852 18228 33908 18284
rect 21746 18172 21756 18228
rect 21812 18172 22540 18228
rect 22596 18172 26908 18228
rect 26964 18172 29036 18228
rect 29092 18172 29102 18228
rect 33842 18172 33852 18228
rect 33908 18172 33918 18228
rect 35186 18172 35196 18228
rect 35252 18172 36932 18228
rect 9650 18060 9660 18116
rect 9716 18060 11676 18116
rect 11732 18060 17892 18116
rect 30930 18060 30940 18116
rect 30996 18060 31006 18116
rect 32162 18060 32172 18116
rect 32228 18060 34636 18116
rect 34692 18060 34702 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 30940 18004 30996 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 14578 17948 14588 18004
rect 14644 17948 15708 18004
rect 15764 17948 16828 18004
rect 16884 17948 16894 18004
rect 19282 17948 19292 18004
rect 19348 17948 20188 18004
rect 20244 17948 21532 18004
rect 21588 17948 21598 18004
rect 26852 17948 33180 18004
rect 33236 17948 33246 18004
rect 20598 17836 20636 17892
rect 20692 17836 20702 17892
rect 24322 17836 24332 17892
rect 24388 17836 24556 17892
rect 24612 17836 24622 17892
rect 11890 17724 11900 17780
rect 11956 17724 13580 17780
rect 13636 17724 13646 17780
rect 14690 17724 14700 17780
rect 14756 17724 23660 17780
rect 23716 17724 23726 17780
rect 26852 17668 26908 17948
rect 36876 17892 36932 18172
rect 36988 18116 37044 18284
rect 38444 18228 38500 18396
rect 39554 18284 39564 18340
rect 39620 18284 41916 18340
rect 41972 18284 42644 18340
rect 42914 18284 42924 18340
rect 42980 18284 44156 18340
rect 44212 18284 44604 18340
rect 44660 18284 44670 18340
rect 42588 18228 42644 18284
rect 38434 18172 38444 18228
rect 38500 18172 38510 18228
rect 42578 18172 42588 18228
rect 42644 18172 42654 18228
rect 36988 18060 37772 18116
rect 37828 18060 39676 18116
rect 39732 18060 39742 18116
rect 30370 17836 30380 17892
rect 30436 17836 30716 17892
rect 30772 17836 31052 17892
rect 31108 17836 36652 17892
rect 36708 17836 36718 17892
rect 36876 17836 42812 17892
rect 42868 17836 43260 17892
rect 43316 17836 43326 17892
rect 28242 17724 28252 17780
rect 28308 17724 31948 17780
rect 32004 17724 32014 17780
rect 33730 17724 33740 17780
rect 33796 17724 34524 17780
rect 34580 17724 34590 17780
rect 36530 17724 36540 17780
rect 36596 17724 37548 17780
rect 37604 17724 37614 17780
rect 38612 17724 41020 17780
rect 41076 17724 41086 17780
rect 38612 17668 38668 17724
rect 7522 17612 7532 17668
rect 7588 17612 7980 17668
rect 8036 17612 8046 17668
rect 10658 17612 10668 17668
rect 10724 17612 15260 17668
rect 15316 17612 15326 17668
rect 15810 17612 15820 17668
rect 15876 17612 17612 17668
rect 17668 17612 17678 17668
rect 17938 17612 17948 17668
rect 18004 17612 18620 17668
rect 18676 17612 18686 17668
rect 18834 17612 18844 17668
rect 18900 17612 23772 17668
rect 23828 17612 23838 17668
rect 24098 17612 24108 17668
rect 24164 17612 25116 17668
rect 25172 17612 25182 17668
rect 26226 17612 26236 17668
rect 26292 17612 26908 17668
rect 27206 17612 27244 17668
rect 27300 17612 27310 17668
rect 30706 17612 30716 17668
rect 30772 17612 31724 17668
rect 31780 17612 33068 17668
rect 33124 17612 33134 17668
rect 35074 17612 35084 17668
rect 35140 17612 38668 17668
rect 38770 17612 38780 17668
rect 38836 17612 39900 17668
rect 39956 17612 39966 17668
rect 45490 17612 45500 17668
rect 45556 17612 47068 17668
rect 47124 17612 47134 17668
rect 59200 17556 60000 17584
rect 13010 17500 13020 17556
rect 13076 17500 14364 17556
rect 14420 17500 14430 17556
rect 16268 17500 23436 17556
rect 23492 17500 24220 17556
rect 24276 17500 24286 17556
rect 30930 17500 30940 17556
rect 30996 17500 31836 17556
rect 31892 17500 31902 17556
rect 33282 17500 33292 17556
rect 33348 17500 34748 17556
rect 34804 17500 34814 17556
rect 41122 17500 41132 17556
rect 41188 17500 41804 17556
rect 41860 17500 41870 17556
rect 42690 17500 42700 17556
rect 42756 17500 45164 17556
rect 45220 17500 45230 17556
rect 57922 17500 57932 17556
rect 57988 17500 60000 17556
rect 16268 17444 16324 17500
rect 59200 17472 60000 17500
rect 7970 17388 7980 17444
rect 8036 17388 8876 17444
rect 8932 17388 8942 17444
rect 13906 17388 13916 17444
rect 13972 17388 14252 17444
rect 14308 17388 14318 17444
rect 14578 17388 14588 17444
rect 14644 17388 16268 17444
rect 16324 17388 16334 17444
rect 18956 17388 21868 17444
rect 21924 17388 21934 17444
rect 24770 17388 24780 17444
rect 24836 17388 26908 17444
rect 26964 17388 26974 17444
rect 27318 17388 27356 17444
rect 27412 17388 27422 17444
rect 27682 17388 27692 17444
rect 27748 17388 27916 17444
rect 27972 17388 27982 17444
rect 28130 17388 28140 17444
rect 28196 17388 29036 17444
rect 29092 17388 29102 17444
rect 32610 17388 32620 17444
rect 32676 17388 32956 17444
rect 33012 17388 33404 17444
rect 33460 17388 33628 17444
rect 33684 17388 33694 17444
rect 39106 17388 39116 17444
rect 39172 17388 39676 17444
rect 39732 17388 41244 17444
rect 41300 17388 41692 17444
rect 41748 17388 41758 17444
rect 42018 17388 42028 17444
rect 42084 17388 46956 17444
rect 47012 17388 47022 17444
rect 47618 17388 47628 17444
rect 47684 17388 47964 17444
rect 48020 17388 48030 17444
rect 18956 17332 19012 17388
rect 10098 17276 10108 17332
rect 10164 17276 15820 17332
rect 15876 17276 15886 17332
rect 17826 17276 17836 17332
rect 17892 17276 18956 17332
rect 19012 17276 19022 17332
rect 20178 17276 20188 17332
rect 20244 17276 20300 17332
rect 20356 17276 22988 17332
rect 23044 17276 23054 17332
rect 23762 17276 23772 17332
rect 23828 17276 35980 17332
rect 36036 17276 37212 17332
rect 37268 17276 37278 17332
rect 38882 17276 38892 17332
rect 38948 17276 41916 17332
rect 41972 17276 41982 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 16482 17164 16492 17220
rect 16548 17164 18844 17220
rect 18900 17164 18910 17220
rect 20738 17164 20748 17220
rect 20804 17164 21196 17220
rect 21252 17164 25228 17220
rect 25284 17164 29596 17220
rect 29652 17164 30268 17220
rect 30324 17164 30334 17220
rect 32050 17164 32060 17220
rect 32116 17164 34188 17220
rect 34244 17164 34254 17220
rect 38658 17164 38668 17220
rect 38724 17164 42812 17220
rect 42868 17164 42878 17220
rect 5394 17052 5404 17108
rect 5460 17052 8428 17108
rect 8484 17052 8494 17108
rect 9874 17052 9884 17108
rect 9940 17052 11900 17108
rect 11956 17052 15036 17108
rect 15092 17052 15102 17108
rect 17714 17052 17724 17108
rect 17780 17052 19852 17108
rect 19908 17052 19918 17108
rect 22530 17052 22540 17108
rect 22596 17052 24780 17108
rect 24836 17052 24846 17108
rect 26114 17052 26124 17108
rect 26180 17052 27244 17108
rect 27300 17052 27310 17108
rect 28924 17052 29372 17108
rect 29428 17052 29932 17108
rect 29988 17052 29998 17108
rect 30482 17052 30492 17108
rect 30548 17052 31052 17108
rect 31108 17052 31118 17108
rect 32386 17052 32396 17108
rect 32452 17052 33404 17108
rect 33460 17052 34300 17108
rect 34356 17052 34366 17108
rect 36866 17052 36876 17108
rect 36932 17052 38108 17108
rect 38164 17052 39788 17108
rect 39844 17052 39854 17108
rect 47058 17052 47068 17108
rect 47124 17052 47964 17108
rect 48020 17052 48030 17108
rect 52098 17052 52108 17108
rect 52164 17052 54460 17108
rect 54516 17052 54526 17108
rect 28924 16996 28980 17052
rect 6402 16940 6412 16996
rect 6468 16940 7644 16996
rect 7700 16940 8316 16996
rect 8372 16940 8382 16996
rect 8978 16940 8988 16996
rect 9044 16940 10500 16996
rect 12002 16940 12012 16996
rect 12068 16940 12348 16996
rect 12404 16940 12414 16996
rect 13794 16940 13804 16996
rect 13860 16940 17388 16996
rect 17444 16940 17454 16996
rect 17724 16940 28980 16996
rect 29138 16940 29148 16996
rect 29204 16940 30156 16996
rect 30212 16940 30828 16996
rect 30884 16940 30894 16996
rect 33170 16940 33180 16996
rect 33236 16940 34412 16996
rect 34468 16940 34478 16996
rect 37986 16940 37996 16996
rect 38052 16940 39116 16996
rect 39172 16940 39182 16996
rect 0 16884 800 16912
rect 10444 16884 10500 16940
rect 0 16828 1708 16884
rect 1764 16828 1774 16884
rect 6066 16828 6076 16884
rect 6132 16828 6972 16884
rect 7028 16828 7038 16884
rect 8306 16828 8316 16884
rect 8372 16828 9324 16884
rect 9380 16828 9390 16884
rect 10434 16828 10444 16884
rect 10500 16828 12516 16884
rect 14578 16828 14588 16884
rect 14644 16828 15484 16884
rect 15540 16828 15550 16884
rect 0 16800 800 16828
rect 12460 16772 12516 16828
rect 17724 16772 17780 16940
rect 18274 16828 18284 16884
rect 18340 16828 20300 16884
rect 20356 16828 20366 16884
rect 23202 16828 23212 16884
rect 23268 16828 25676 16884
rect 25732 16828 25742 16884
rect 27122 16828 27132 16884
rect 27188 16828 27804 16884
rect 27860 16828 27870 16884
rect 28588 16828 31500 16884
rect 31556 16828 31566 16884
rect 37538 16828 37548 16884
rect 37604 16828 37772 16884
rect 37828 16828 41468 16884
rect 41524 16828 42140 16884
rect 42196 16828 42206 16884
rect 51538 16828 51548 16884
rect 51604 16828 53340 16884
rect 53396 16828 54572 16884
rect 54628 16828 54638 16884
rect 28588 16772 28644 16828
rect 7298 16716 7308 16772
rect 7364 16716 8428 16772
rect 8484 16716 8494 16772
rect 12450 16716 12460 16772
rect 12516 16716 13468 16772
rect 13524 16716 13804 16772
rect 13860 16716 13870 16772
rect 14130 16716 14140 16772
rect 14196 16716 17780 16772
rect 22194 16716 22204 16772
rect 22260 16716 22540 16772
rect 22596 16716 22606 16772
rect 23538 16716 23548 16772
rect 23604 16716 23884 16772
rect 23940 16716 26460 16772
rect 26516 16716 26526 16772
rect 27570 16716 27580 16772
rect 27636 16716 28644 16772
rect 34374 16716 34412 16772
rect 34468 16716 34478 16772
rect 35298 16716 35308 16772
rect 35364 16716 38668 16772
rect 38882 16716 38892 16772
rect 38948 16716 40124 16772
rect 40180 16716 40190 16772
rect 40338 16716 40348 16772
rect 40404 16716 41356 16772
rect 41412 16716 41422 16772
rect 41794 16716 41804 16772
rect 41860 16716 45052 16772
rect 45108 16716 45118 16772
rect 45490 16716 45500 16772
rect 45556 16716 46060 16772
rect 46116 16716 46126 16772
rect 38612 16660 38668 16716
rect 10098 16604 10108 16660
rect 10164 16604 16156 16660
rect 16212 16604 19180 16660
rect 19236 16604 19246 16660
rect 24098 16604 24108 16660
rect 24164 16604 29372 16660
rect 29428 16604 29438 16660
rect 34850 16604 34860 16660
rect 34916 16604 35196 16660
rect 35252 16604 35262 16660
rect 38612 16604 40908 16660
rect 40964 16604 40974 16660
rect 41356 16548 41412 16716
rect 41906 16604 41916 16660
rect 41972 16604 48188 16660
rect 48244 16604 48254 16660
rect 52770 16604 52780 16660
rect 52836 16604 54236 16660
rect 54292 16604 54302 16660
rect 5842 16492 5852 16548
rect 5908 16492 10332 16548
rect 10388 16492 13468 16548
rect 13524 16492 14140 16548
rect 14196 16492 14206 16548
rect 15586 16492 15596 16548
rect 15652 16492 17164 16548
rect 17220 16492 20580 16548
rect 22978 16492 22988 16548
rect 23044 16492 25004 16548
rect 25060 16492 25070 16548
rect 27346 16492 27356 16548
rect 27412 16492 29148 16548
rect 29204 16492 29214 16548
rect 41356 16492 42028 16548
rect 42084 16492 42364 16548
rect 42420 16492 42430 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 20524 16436 20580 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 12898 16380 12908 16436
rect 12964 16380 18172 16436
rect 18228 16380 20188 16436
rect 20244 16380 20254 16436
rect 20514 16380 20524 16436
rect 20580 16380 20860 16436
rect 20916 16380 20926 16436
rect 24322 16380 24332 16436
rect 24388 16380 25676 16436
rect 25732 16380 25742 16436
rect 32918 16380 32956 16436
rect 33012 16380 33516 16436
rect 33572 16380 33740 16436
rect 33796 16380 33806 16436
rect 8194 16268 8204 16324
rect 8260 16268 10780 16324
rect 10836 16268 10846 16324
rect 15362 16268 15372 16324
rect 15428 16268 17276 16324
rect 17332 16268 17342 16324
rect 20066 16268 20076 16324
rect 20132 16268 20972 16324
rect 21028 16268 26908 16324
rect 26964 16268 26974 16324
rect 27542 16268 27580 16324
rect 27636 16268 27646 16324
rect 28914 16268 28924 16324
rect 28980 16268 29484 16324
rect 29540 16268 29550 16324
rect 31826 16268 31836 16324
rect 31892 16268 40348 16324
rect 40404 16268 40414 16324
rect 12002 16156 12012 16212
rect 12068 16156 13356 16212
rect 13412 16156 15372 16212
rect 15428 16156 16716 16212
rect 16772 16156 16782 16212
rect 17378 16156 17388 16212
rect 17444 16156 18172 16212
rect 18228 16156 22652 16212
rect 22708 16156 22718 16212
rect 26562 16156 26572 16212
rect 26628 16156 39564 16212
rect 39620 16156 39630 16212
rect 42466 16156 42476 16212
rect 42532 16156 49532 16212
rect 49588 16156 50092 16212
rect 50148 16156 50158 16212
rect 50978 16156 50988 16212
rect 51044 16156 51772 16212
rect 51828 16156 53004 16212
rect 53060 16156 53070 16212
rect 14802 16044 14812 16100
rect 14868 16044 15148 16100
rect 15204 16044 15214 16100
rect 15810 16044 15820 16100
rect 15876 16044 19964 16100
rect 20020 16044 20030 16100
rect 22754 16044 22764 16100
rect 22820 16044 23212 16100
rect 23268 16044 23278 16100
rect 25330 16044 25340 16100
rect 25396 16044 25788 16100
rect 25844 16044 25854 16100
rect 26674 16044 26684 16100
rect 26740 16044 27468 16100
rect 27524 16044 27534 16100
rect 31826 16044 31836 16100
rect 31892 16044 33404 16100
rect 33460 16044 33470 16100
rect 43026 16044 43036 16100
rect 43092 16044 43596 16100
rect 43652 16044 43932 16100
rect 43988 16044 43998 16100
rect 44146 16044 44156 16100
rect 44212 16044 46172 16100
rect 46228 16044 46238 16100
rect 47170 16044 47180 16100
rect 47236 16044 47516 16100
rect 47572 16044 47582 16100
rect 51538 16044 51548 16100
rect 51604 16044 52892 16100
rect 52948 16044 52958 16100
rect 5730 15932 5740 15988
rect 5796 15932 6524 15988
rect 6580 15932 6972 15988
rect 7028 15932 7038 15988
rect 11218 15932 11228 15988
rect 11284 15932 11676 15988
rect 11732 15932 11742 15988
rect 15026 15932 15036 15988
rect 15092 15932 16660 15988
rect 18834 15932 18844 15988
rect 18900 15932 22092 15988
rect 22148 15932 22158 15988
rect 23090 15932 23100 15988
rect 23156 15932 24780 15988
rect 24836 15932 24846 15988
rect 26450 15932 26460 15988
rect 26516 15932 28812 15988
rect 28868 15932 32060 15988
rect 32116 15932 32126 15988
rect 43362 15932 43372 15988
rect 43428 15932 44828 15988
rect 44884 15932 44894 15988
rect 16604 15876 16660 15932
rect 11106 15820 11116 15876
rect 11172 15820 15652 15876
rect 15810 15820 15820 15876
rect 15876 15820 16156 15876
rect 16212 15820 16222 15876
rect 16594 15820 16604 15876
rect 16660 15820 17948 15876
rect 18004 15820 18284 15876
rect 18340 15820 18350 15876
rect 19618 15820 19628 15876
rect 19684 15820 21308 15876
rect 21364 15820 21374 15876
rect 22306 15820 22316 15876
rect 22372 15820 23436 15876
rect 23492 15820 27356 15876
rect 27412 15820 27422 15876
rect 28130 15820 28140 15876
rect 28196 15820 37100 15876
rect 37156 15820 37436 15876
rect 37492 15820 37884 15876
rect 37940 15820 38220 15876
rect 38276 15820 38668 15876
rect 42690 15820 42700 15876
rect 42756 15820 46732 15876
rect 46788 15820 47068 15876
rect 47124 15820 47134 15876
rect 48066 15820 48076 15876
rect 48132 15820 49084 15876
rect 49140 15820 49150 15876
rect 49634 15820 49644 15876
rect 49700 15820 51212 15876
rect 51268 15820 51278 15876
rect 15596 15764 15652 15820
rect 10434 15708 10444 15764
rect 10500 15708 15372 15764
rect 15428 15708 15438 15764
rect 15596 15708 16268 15764
rect 16324 15708 16334 15764
rect 22530 15708 22540 15764
rect 22596 15708 25620 15764
rect 28578 15708 28588 15764
rect 28644 15708 29932 15764
rect 29988 15708 31164 15764
rect 31220 15708 31230 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 25564 15652 25620 15708
rect 38612 15652 38668 15820
rect 45154 15708 45164 15764
rect 45220 15708 46508 15764
rect 46564 15708 46574 15764
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 13682 15596 13692 15652
rect 13748 15596 14812 15652
rect 14868 15596 14878 15652
rect 15362 15596 15372 15652
rect 15428 15596 18508 15652
rect 18564 15596 18574 15652
rect 22306 15596 22316 15652
rect 22372 15596 22652 15652
rect 22708 15596 22718 15652
rect 25564 15596 25676 15652
rect 25732 15596 26460 15652
rect 26516 15596 26526 15652
rect 26852 15596 35868 15652
rect 35924 15596 36988 15652
rect 37044 15596 37054 15652
rect 37426 15596 37436 15652
rect 37492 15596 38108 15652
rect 38164 15596 38174 15652
rect 38612 15596 38892 15652
rect 38948 15596 38958 15652
rect 26852 15540 26908 15596
rect 14578 15484 14588 15540
rect 14644 15484 15596 15540
rect 15652 15484 15662 15540
rect 16706 15484 16716 15540
rect 16772 15484 26908 15540
rect 27346 15484 27356 15540
rect 27412 15484 30380 15540
rect 30436 15484 32396 15540
rect 32452 15484 32462 15540
rect 37090 15484 37100 15540
rect 37156 15484 38332 15540
rect 38388 15484 38398 15540
rect 7746 15372 7756 15428
rect 7812 15372 9548 15428
rect 9604 15372 9614 15428
rect 10098 15372 10108 15428
rect 10164 15372 11788 15428
rect 11844 15372 11854 15428
rect 12012 15372 15036 15428
rect 15092 15372 15102 15428
rect 16258 15372 16268 15428
rect 16324 15372 18956 15428
rect 19012 15372 23100 15428
rect 23156 15372 23166 15428
rect 28242 15372 28252 15428
rect 28308 15372 28588 15428
rect 28644 15372 30156 15428
rect 30212 15372 30222 15428
rect 33730 15372 33740 15428
rect 33796 15372 34076 15428
rect 34132 15372 34142 15428
rect 36866 15372 36876 15428
rect 36932 15372 37324 15428
rect 37380 15372 37390 15428
rect 42018 15372 42028 15428
rect 42084 15372 42476 15428
rect 42532 15372 42542 15428
rect 52658 15372 52668 15428
rect 52724 15372 53564 15428
rect 53620 15372 53630 15428
rect 12012 15316 12068 15372
rect 5618 15260 5628 15316
rect 5684 15260 7084 15316
rect 7140 15260 12068 15316
rect 12124 15260 16604 15316
rect 16660 15260 16772 15316
rect 17266 15260 17276 15316
rect 17332 15260 19964 15316
rect 20020 15260 20030 15316
rect 21410 15260 21420 15316
rect 21476 15260 22764 15316
rect 22820 15260 22830 15316
rect 24294 15260 24332 15316
rect 24388 15260 24398 15316
rect 25788 15260 26124 15316
rect 26180 15260 27692 15316
rect 27748 15260 27758 15316
rect 28662 15260 28700 15316
rect 28756 15260 28766 15316
rect 32162 15260 32172 15316
rect 32228 15260 33180 15316
rect 33236 15260 33246 15316
rect 33618 15260 33628 15316
rect 33684 15260 34636 15316
rect 34692 15260 34702 15316
rect 41458 15260 41468 15316
rect 41524 15260 42924 15316
rect 42980 15260 42990 15316
rect 49410 15260 49420 15316
rect 49476 15260 50988 15316
rect 51044 15260 51054 15316
rect 12124 15204 12180 15260
rect 8418 15148 8428 15204
rect 8484 15148 12180 15204
rect 15026 15148 15036 15204
rect 15092 15148 15820 15204
rect 15876 15148 15886 15204
rect 16716 15092 16772 15260
rect 19964 15204 20020 15260
rect 25788 15204 25844 15260
rect 19964 15148 25788 15204
rect 25844 15148 25854 15204
rect 36978 15148 36988 15204
rect 37044 15148 38556 15204
rect 38612 15148 41244 15204
rect 41300 15148 41310 15204
rect 49074 15148 49084 15204
rect 49140 15148 49980 15204
rect 50036 15148 50046 15204
rect 41244 15092 41300 15148
rect 7970 15036 7980 15092
rect 8036 15036 8204 15092
rect 8260 15036 8270 15092
rect 9986 15036 9996 15092
rect 10052 15036 11788 15092
rect 11844 15036 12796 15092
rect 12852 15036 13804 15092
rect 13860 15036 13870 15092
rect 14466 15036 14476 15092
rect 14532 15036 16492 15092
rect 16548 15036 16558 15092
rect 16716 15036 17108 15092
rect 18722 15036 18732 15092
rect 18788 15036 19404 15092
rect 19460 15036 19470 15092
rect 19842 15036 19852 15092
rect 19908 15036 26572 15092
rect 26628 15036 27804 15092
rect 27860 15036 27870 15092
rect 34402 15036 34412 15092
rect 34468 15036 34972 15092
rect 35028 15036 35038 15092
rect 37090 15036 37100 15092
rect 37156 15036 37660 15092
rect 37716 15036 37726 15092
rect 41244 15036 42028 15092
rect 42084 15036 42094 15092
rect 48850 15036 48860 15092
rect 48916 15036 49756 15092
rect 49812 15036 49822 15092
rect 17052 14980 17108 15036
rect 8306 14924 8316 14980
rect 8372 14924 12908 14980
rect 12964 14924 16044 14980
rect 16100 14924 16110 14980
rect 17052 14924 17388 14980
rect 17444 14924 27580 14980
rect 27636 14924 28588 14980
rect 28644 14924 28700 14980
rect 28756 14924 30156 14980
rect 30212 14924 31836 14980
rect 31892 14924 31902 14980
rect 33478 14924 33516 14980
rect 33572 14924 33582 14980
rect 37538 14924 37548 14980
rect 37604 14924 38108 14980
rect 38164 14924 38174 14980
rect 39330 14924 39340 14980
rect 39396 14924 40236 14980
rect 40292 14924 40302 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 59200 14868 60000 14896
rect 6850 14812 6860 14868
rect 6916 14812 7868 14868
rect 7924 14812 7934 14868
rect 11330 14812 11340 14868
rect 11396 14812 20188 14868
rect 20244 14812 21532 14868
rect 21588 14812 21598 14868
rect 31052 14812 35028 14868
rect 39778 14812 39788 14868
rect 39844 14812 41020 14868
rect 41076 14812 41086 14868
rect 45938 14812 45948 14868
rect 46004 14812 46014 14868
rect 46470 14812 46508 14868
rect 46564 14812 46574 14868
rect 57922 14812 57932 14868
rect 57988 14812 60000 14868
rect 31052 14756 31108 14812
rect 34972 14756 35028 14812
rect 6290 14700 6300 14756
rect 6356 14700 7644 14756
rect 7700 14700 7710 14756
rect 9090 14700 9100 14756
rect 9156 14700 10108 14756
rect 10164 14700 10668 14756
rect 10724 14700 10734 14756
rect 17154 14700 17164 14756
rect 17220 14700 18396 14756
rect 18452 14700 18462 14756
rect 18722 14700 18732 14756
rect 18788 14700 19852 14756
rect 19908 14700 19918 14756
rect 21298 14700 21308 14756
rect 21364 14700 31108 14756
rect 31266 14700 31276 14756
rect 31332 14700 31836 14756
rect 31892 14700 31902 14756
rect 34972 14700 36428 14756
rect 36484 14700 36494 14756
rect 38658 14700 38668 14756
rect 38724 14700 39900 14756
rect 39956 14700 39966 14756
rect 17164 14644 17220 14700
rect 6738 14588 6748 14644
rect 6804 14588 9548 14644
rect 9604 14588 13468 14644
rect 13524 14588 13534 14644
rect 15362 14588 15372 14644
rect 15428 14588 17220 14644
rect 18162 14588 18172 14644
rect 18228 14588 19292 14644
rect 19348 14588 24668 14644
rect 24724 14588 27356 14644
rect 27412 14588 27422 14644
rect 29810 14588 29820 14644
rect 29876 14588 31388 14644
rect 31444 14588 31948 14644
rect 32004 14588 32014 14644
rect 6178 14476 6188 14532
rect 6244 14476 9212 14532
rect 9268 14476 10332 14532
rect 10388 14476 10398 14532
rect 14914 14476 14924 14532
rect 14980 14476 15932 14532
rect 15988 14476 15998 14532
rect 22978 14476 22988 14532
rect 23044 14476 23324 14532
rect 23380 14476 23436 14532
rect 23492 14476 25172 14532
rect 25666 14476 25676 14532
rect 25732 14476 27468 14532
rect 27524 14476 27534 14532
rect 28242 14476 28252 14532
rect 28308 14476 28318 14532
rect 28466 14476 28476 14532
rect 28532 14476 31276 14532
rect 31332 14476 31342 14532
rect 36418 14476 36428 14532
rect 36484 14476 45500 14532
rect 45556 14476 45566 14532
rect 25116 14420 25172 14476
rect 28252 14420 28308 14476
rect 45948 14420 46004 14812
rect 59200 14784 60000 14812
rect 54562 14476 54572 14532
rect 54628 14476 55580 14532
rect 55636 14476 55646 14532
rect 9762 14364 9772 14420
rect 9828 14364 10444 14420
rect 10500 14364 11228 14420
rect 11284 14364 11294 14420
rect 13682 14364 13692 14420
rect 13748 14364 24444 14420
rect 24500 14364 24892 14420
rect 24948 14364 24958 14420
rect 25116 14364 27132 14420
rect 27188 14364 27198 14420
rect 27682 14364 27692 14420
rect 27748 14364 28308 14420
rect 29698 14364 29708 14420
rect 29764 14364 31724 14420
rect 31780 14364 31790 14420
rect 32946 14364 32956 14420
rect 33012 14364 34188 14420
rect 34244 14364 34254 14420
rect 37090 14364 37100 14420
rect 37156 14364 37660 14420
rect 37716 14364 37726 14420
rect 38434 14364 38444 14420
rect 38500 14364 40124 14420
rect 40180 14364 40190 14420
rect 43138 14364 43148 14420
rect 43204 14364 46732 14420
rect 46788 14364 46798 14420
rect 50866 14364 50876 14420
rect 50932 14364 51660 14420
rect 51716 14364 52220 14420
rect 52276 14364 52286 14420
rect 38444 14308 38500 14364
rect 9874 14252 9884 14308
rect 9940 14252 13804 14308
rect 13860 14252 14476 14308
rect 14532 14252 14542 14308
rect 19628 14252 19740 14308
rect 19796 14252 19806 14308
rect 23426 14252 23436 14308
rect 23492 14252 26012 14308
rect 26068 14252 29148 14308
rect 29204 14252 29214 14308
rect 34738 14252 34748 14308
rect 34804 14252 35420 14308
rect 35476 14252 35486 14308
rect 36642 14252 36652 14308
rect 36708 14252 37884 14308
rect 37940 14252 38500 14308
rect 42802 14252 42812 14308
rect 42868 14252 43484 14308
rect 43540 14252 43550 14308
rect 46470 14252 46508 14308
rect 46564 14252 46574 14308
rect 19628 14196 19684 14252
rect 10210 14140 10220 14196
rect 10276 14140 10668 14196
rect 10724 14140 11900 14196
rect 11956 14140 12684 14196
rect 12740 14140 13244 14196
rect 13300 14140 13310 14196
rect 19618 14140 19628 14196
rect 19684 14140 19694 14196
rect 27878 14140 27916 14196
rect 27972 14140 27982 14196
rect 28914 14140 28924 14196
rect 28980 14140 31612 14196
rect 31668 14140 34972 14196
rect 35028 14140 36428 14196
rect 36484 14140 36494 14196
rect 46246 14140 46284 14196
rect 46340 14140 46350 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 6962 14028 6972 14084
rect 7028 14028 8204 14084
rect 8260 14028 15372 14084
rect 15428 14028 15438 14084
rect 17126 14028 17164 14084
rect 17220 14028 17230 14084
rect 27682 14028 27692 14084
rect 27748 14028 29372 14084
rect 29428 14028 29438 14084
rect 38322 14028 38332 14084
rect 38388 14028 40012 14084
rect 40068 14028 40078 14084
rect 8530 13916 8540 13972
rect 8596 13916 8606 13972
rect 13010 13916 13020 13972
rect 13076 13916 14588 13972
rect 14644 13916 14654 13972
rect 15586 13916 15596 13972
rect 15652 13916 16044 13972
rect 16100 13916 16110 13972
rect 18386 13916 18396 13972
rect 18452 13916 20132 13972
rect 23538 13916 23548 13972
rect 23604 13916 23772 13972
rect 23828 13916 23838 13972
rect 24658 13916 24668 13972
rect 24724 13916 28028 13972
rect 28084 13916 28094 13972
rect 8540 13748 8596 13916
rect 20076 13860 20132 13916
rect 12786 13804 12796 13860
rect 12852 13804 19852 13860
rect 19908 13804 19918 13860
rect 20076 13804 25452 13860
rect 25508 13804 25518 13860
rect 25778 13804 25788 13860
rect 25844 13804 34076 13860
rect 34132 13804 34142 13860
rect 46050 13804 46060 13860
rect 46116 13804 47180 13860
rect 47236 13804 47246 13860
rect 7186 13692 7196 13748
rect 7252 13692 8092 13748
rect 8148 13692 8158 13748
rect 8540 13692 9772 13748
rect 9828 13692 9838 13748
rect 10434 13692 10444 13748
rect 10500 13692 10668 13748
rect 10724 13692 11452 13748
rect 11508 13692 11518 13748
rect 14018 13692 14028 13748
rect 14084 13692 14700 13748
rect 14756 13692 14766 13748
rect 16818 13692 16828 13748
rect 16884 13692 18060 13748
rect 18116 13692 18126 13748
rect 27346 13692 27356 13748
rect 27412 13692 31052 13748
rect 31108 13692 31118 13748
rect 32498 13692 32508 13748
rect 32564 13692 35532 13748
rect 35588 13692 35598 13748
rect 37548 13692 38668 13748
rect 38724 13692 38734 13748
rect 39890 13692 39900 13748
rect 39956 13692 45388 13748
rect 45444 13692 45454 13748
rect 6514 13580 6524 13636
rect 6580 13580 7644 13636
rect 7700 13580 8204 13636
rect 8260 13580 8270 13636
rect 18134 13580 18172 13636
rect 18228 13580 18238 13636
rect 19394 13580 19404 13636
rect 19460 13580 21196 13636
rect 21252 13580 21262 13636
rect 30818 13580 30828 13636
rect 30884 13580 31724 13636
rect 31780 13580 31790 13636
rect 32274 13580 32284 13636
rect 32340 13580 32732 13636
rect 32788 13580 33180 13636
rect 33236 13580 33246 13636
rect 35074 13580 35084 13636
rect 35140 13580 37100 13636
rect 37156 13580 37166 13636
rect 37548 13524 37604 13692
rect 40898 13580 40908 13636
rect 40964 13580 42924 13636
rect 42980 13580 42990 13636
rect 5954 13468 5964 13524
rect 6020 13468 7028 13524
rect 7186 13468 7196 13524
rect 7252 13468 8540 13524
rect 8596 13468 8606 13524
rect 14914 13468 14924 13524
rect 14980 13468 15260 13524
rect 15316 13468 15326 13524
rect 15474 13468 15484 13524
rect 15540 13468 16884 13524
rect 25218 13468 25228 13524
rect 25284 13468 28476 13524
rect 28532 13468 28542 13524
rect 31042 13468 31052 13524
rect 31108 13468 33852 13524
rect 33908 13468 33918 13524
rect 37538 13468 37548 13524
rect 37604 13468 37614 13524
rect 37762 13468 37772 13524
rect 37828 13468 38892 13524
rect 38948 13468 41020 13524
rect 41076 13468 41086 13524
rect 42018 13468 42028 13524
rect 42084 13468 42812 13524
rect 42868 13468 42878 13524
rect 6972 13412 7028 13468
rect 16828 13412 16884 13468
rect 6972 13356 7084 13412
rect 7140 13356 7150 13412
rect 7522 13356 7532 13412
rect 7588 13356 8876 13412
rect 8932 13356 8942 13412
rect 16828 13356 18732 13412
rect 18788 13356 18798 13412
rect 22642 13356 22652 13412
rect 22708 13356 23324 13412
rect 23380 13356 23390 13412
rect 25106 13356 25116 13412
rect 25172 13356 33404 13412
rect 33460 13356 33470 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 22754 13244 22764 13300
rect 22820 13244 24108 13300
rect 24164 13244 24174 13300
rect 25554 13244 25564 13300
rect 25620 13244 26124 13300
rect 26180 13244 26190 13300
rect 28242 13244 28252 13300
rect 28308 13244 33628 13300
rect 33684 13244 33694 13300
rect 11554 13132 11564 13188
rect 11620 13132 34300 13188
rect 34356 13132 37548 13188
rect 37604 13132 37614 13188
rect 6738 13020 6748 13076
rect 6804 13020 12012 13076
rect 12068 13020 12078 13076
rect 14214 13020 14252 13076
rect 14308 13020 14318 13076
rect 14466 13020 14476 13076
rect 14532 13020 14570 13076
rect 19842 13020 19852 13076
rect 19908 13020 21196 13076
rect 21252 13020 21262 13076
rect 24994 13020 25004 13076
rect 25060 13020 28252 13076
rect 28308 13020 28318 13076
rect 30258 13020 30268 13076
rect 30324 13020 31948 13076
rect 32004 13020 32014 13076
rect 38434 13020 38444 13076
rect 38500 13020 38510 13076
rect 40674 13020 40684 13076
rect 40740 13020 42364 13076
rect 42420 13020 42430 13076
rect 51650 13020 51660 13076
rect 51716 13020 52780 13076
rect 52836 13020 52846 13076
rect 6290 12908 6300 12964
rect 6356 12908 6636 12964
rect 6692 12908 7084 12964
rect 7140 12908 7150 12964
rect 14354 12908 14364 12964
rect 14420 12908 15036 12964
rect 15092 12908 15102 12964
rect 16258 12908 16268 12964
rect 16324 12908 16940 12964
rect 16996 12908 17006 12964
rect 20626 12908 20636 12964
rect 20692 12908 21868 12964
rect 21924 12908 23436 12964
rect 23492 12908 23502 12964
rect 26114 12908 26124 12964
rect 26180 12908 26908 12964
rect 26964 12908 26974 12964
rect 30706 12908 30716 12964
rect 30772 12908 31388 12964
rect 31444 12908 35644 12964
rect 35700 12908 35710 12964
rect 37650 12908 37660 12964
rect 37716 12908 38220 12964
rect 38276 12908 38286 12964
rect 38444 12852 38500 13020
rect 40450 12908 40460 12964
rect 40516 12908 43372 12964
rect 43428 12908 43932 12964
rect 43988 12908 44268 12964
rect 44324 12908 44334 12964
rect 51314 12908 51324 12964
rect 51380 12908 53004 12964
rect 53060 12908 53070 12964
rect 7410 12796 7420 12852
rect 7476 12796 8428 12852
rect 8484 12796 8494 12852
rect 9650 12796 9660 12852
rect 9716 12796 10108 12852
rect 10164 12796 10174 12852
rect 15092 12796 23324 12852
rect 23380 12796 23772 12852
rect 23828 12796 23838 12852
rect 25442 12796 25452 12852
rect 25508 12796 27188 12852
rect 15092 12740 15148 12796
rect 27132 12740 27188 12796
rect 33740 12796 37100 12852
rect 37156 12796 37166 12852
rect 38220 12796 38500 12852
rect 38612 12796 40012 12852
rect 40068 12796 41468 12852
rect 41524 12796 41534 12852
rect 49746 12796 49756 12852
rect 49812 12796 51100 12852
rect 51156 12796 51772 12852
rect 51828 12796 51838 12852
rect 33740 12740 33796 12796
rect 38220 12740 38276 12796
rect 12338 12684 12348 12740
rect 12404 12684 14588 12740
rect 14644 12684 15148 12740
rect 19058 12684 19068 12740
rect 19124 12684 20188 12740
rect 20244 12684 26908 12740
rect 27122 12684 27132 12740
rect 27188 12684 27198 12740
rect 27906 12684 27916 12740
rect 27972 12684 28028 12740
rect 28084 12684 28094 12740
rect 31378 12684 31388 12740
rect 31444 12684 31454 12740
rect 32722 12684 32732 12740
rect 32788 12684 33516 12740
rect 33572 12684 33796 12740
rect 33954 12684 33964 12740
rect 34020 12684 36316 12740
rect 36372 12684 36382 12740
rect 38210 12684 38220 12740
rect 38276 12684 38286 12740
rect 38546 12684 38556 12740
rect 38612 12684 38668 12796
rect 39442 12684 39452 12740
rect 39508 12684 40124 12740
rect 40180 12684 41692 12740
rect 41748 12684 41758 12740
rect 50978 12684 50988 12740
rect 51044 12684 52108 12740
rect 52164 12684 52174 12740
rect 11106 12572 11116 12628
rect 11172 12572 11452 12628
rect 11508 12572 11518 12628
rect 12226 12572 12236 12628
rect 12292 12572 15148 12628
rect 20486 12572 20524 12628
rect 20580 12572 20590 12628
rect 15092 12516 15148 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 26852 12516 26908 12684
rect 31388 12516 31444 12684
rect 40786 12572 40796 12628
rect 40852 12572 47404 12628
rect 47460 12572 47470 12628
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 8418 12460 8428 12516
rect 8484 12460 13580 12516
rect 13636 12460 13646 12516
rect 15092 12460 19068 12516
rect 19124 12460 19134 12516
rect 26852 12460 27804 12516
rect 27860 12460 27870 12516
rect 31388 12460 41244 12516
rect 41300 12460 42476 12516
rect 42532 12460 42542 12516
rect 9090 12348 9100 12404
rect 9156 12348 12236 12404
rect 12292 12348 12302 12404
rect 12562 12348 12572 12404
rect 12628 12348 17612 12404
rect 17668 12348 17678 12404
rect 18274 12348 18284 12404
rect 18340 12348 38220 12404
rect 38276 12348 39900 12404
rect 39956 12348 39966 12404
rect 45948 12348 48748 12404
rect 48804 12348 48814 12404
rect 49308 12348 50204 12404
rect 50260 12348 50270 12404
rect 51874 12348 51884 12404
rect 51940 12348 52668 12404
rect 52724 12348 52734 12404
rect 45948 12292 46004 12348
rect 49308 12292 49364 12348
rect 10882 12236 10892 12292
rect 10948 12236 12124 12292
rect 12180 12236 12190 12292
rect 15586 12236 15596 12292
rect 15652 12236 16268 12292
rect 16324 12236 19628 12292
rect 19684 12236 19852 12292
rect 19908 12236 19918 12292
rect 20524 12236 21420 12292
rect 21476 12236 22652 12292
rect 22708 12236 22718 12292
rect 28578 12236 28588 12292
rect 28644 12236 31388 12292
rect 31444 12236 31724 12292
rect 31780 12236 31790 12292
rect 37314 12236 37324 12292
rect 37380 12236 46004 12292
rect 46162 12236 46172 12292
rect 46228 12236 48972 12292
rect 49028 12236 49308 12292
rect 49364 12236 49374 12292
rect 49970 12236 49980 12292
rect 50036 12236 50988 12292
rect 51044 12236 51054 12292
rect 7942 12124 7980 12180
rect 8036 12124 8046 12180
rect 11106 12124 11116 12180
rect 11172 12124 12684 12180
rect 12740 12124 19180 12180
rect 19236 12124 19246 12180
rect 20524 12068 20580 12236
rect 59200 12180 60000 12208
rect 20738 12124 20748 12180
rect 20804 12124 20814 12180
rect 22082 12124 22092 12180
rect 22148 12124 22540 12180
rect 22596 12124 22606 12180
rect 23874 12124 23884 12180
rect 23940 12124 29820 12180
rect 29876 12124 29886 12180
rect 34626 12124 34636 12180
rect 34692 12124 35084 12180
rect 35140 12124 35150 12180
rect 35858 12124 35868 12180
rect 35924 12124 36428 12180
rect 36484 12124 36494 12180
rect 39554 12124 39564 12180
rect 39620 12124 40684 12180
rect 40740 12124 40750 12180
rect 43810 12124 43820 12180
rect 43876 12124 45388 12180
rect 45444 12124 45454 12180
rect 48178 12124 48188 12180
rect 48244 12124 48860 12180
rect 48916 12124 49532 12180
rect 49588 12124 50764 12180
rect 50820 12124 50830 12180
rect 52322 12124 52332 12180
rect 52388 12124 53452 12180
rect 53508 12124 53518 12180
rect 53890 12124 53900 12180
rect 53956 12124 54572 12180
rect 54628 12124 54638 12180
rect 57922 12124 57932 12180
rect 57988 12124 60000 12180
rect 6850 12012 6860 12068
rect 6916 12012 11564 12068
rect 11620 12012 11630 12068
rect 12002 12012 12012 12068
rect 12068 12012 20580 12068
rect 20748 11956 20804 12124
rect 59200 12096 60000 12124
rect 22306 12012 22316 12068
rect 22372 12012 23212 12068
rect 23268 12012 23278 12068
rect 28242 12012 28252 12068
rect 28308 12012 29708 12068
rect 29764 12012 29774 12068
rect 42354 12012 42364 12068
rect 42420 12012 42812 12068
rect 42868 12012 42878 12068
rect 8306 11900 8316 11956
rect 8372 11900 20804 11956
rect 21970 11900 21980 11956
rect 22036 11900 25676 11956
rect 25732 11900 25742 11956
rect 28354 11900 28364 11956
rect 28420 11900 35868 11956
rect 35924 11900 35934 11956
rect 42242 11900 42252 11956
rect 42308 11900 43148 11956
rect 43204 11900 43214 11956
rect 8978 11788 8988 11844
rect 9044 11788 10332 11844
rect 10388 11788 12012 11844
rect 12068 11788 12078 11844
rect 14018 11788 14028 11844
rect 14084 11788 16828 11844
rect 16884 11788 16894 11844
rect 20066 11788 20076 11844
rect 20132 11788 20412 11844
rect 20468 11788 20478 11844
rect 20598 11788 20636 11844
rect 20692 11788 20702 11844
rect 21858 11788 21868 11844
rect 21924 11788 25004 11844
rect 25060 11788 25070 11844
rect 34822 11788 34860 11844
rect 34916 11788 34926 11844
rect 47506 11788 47516 11844
rect 47572 11788 48412 11844
rect 48468 11788 48478 11844
rect 54338 11788 54348 11844
rect 54404 11788 55692 11844
rect 55748 11788 55758 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 10780 11676 10892 11732
rect 10948 11676 10958 11732
rect 11442 11676 11452 11732
rect 11508 11676 12572 11732
rect 12628 11676 12638 11732
rect 14578 11676 14588 11732
rect 14644 11676 14924 11732
rect 14980 11676 14990 11732
rect 16706 11676 16716 11732
rect 16772 11676 17836 11732
rect 17892 11676 17902 11732
rect 18162 11676 18172 11732
rect 18228 11676 18956 11732
rect 19012 11676 19022 11732
rect 26114 11676 26124 11732
rect 26180 11676 28364 11732
rect 28420 11676 28430 11732
rect 28578 11676 28588 11732
rect 28644 11676 29820 11732
rect 29876 11676 29886 11732
rect 37762 11676 37772 11732
rect 37828 11676 38780 11732
rect 38836 11676 38846 11732
rect 52098 11676 52108 11732
rect 52164 11676 52780 11732
rect 52836 11676 53788 11732
rect 53844 11676 53854 11732
rect 10780 11620 10836 11676
rect 16716 11620 16772 11676
rect 10658 11564 10668 11620
rect 10724 11564 10836 11620
rect 11218 11564 11228 11620
rect 11284 11564 13692 11620
rect 13748 11564 16772 11620
rect 25106 11564 25116 11620
rect 25172 11564 27860 11620
rect 28690 11564 28700 11620
rect 28756 11564 32172 11620
rect 32228 11564 32238 11620
rect 34514 11564 34524 11620
rect 34580 11564 34972 11620
rect 35028 11564 35038 11620
rect 27804 11508 27860 11564
rect 7522 11452 7532 11508
rect 7588 11452 8764 11508
rect 8820 11452 10108 11508
rect 10164 11452 10780 11508
rect 10836 11452 10846 11508
rect 11452 11452 16940 11508
rect 16996 11452 17006 11508
rect 19030 11452 19068 11508
rect 19124 11452 19134 11508
rect 19282 11452 19292 11508
rect 19348 11452 19852 11508
rect 19908 11452 19918 11508
rect 21634 11452 21644 11508
rect 21700 11452 27580 11508
rect 27636 11452 27646 11508
rect 27804 11452 36092 11508
rect 36148 11452 36158 11508
rect 36866 11452 36876 11508
rect 36932 11452 38444 11508
rect 38500 11452 38510 11508
rect 43250 11452 43260 11508
rect 43316 11452 43484 11508
rect 43540 11452 43550 11508
rect 45154 11452 45164 11508
rect 45220 11452 45724 11508
rect 45780 11452 46396 11508
rect 46452 11452 46462 11508
rect 10322 11340 10332 11396
rect 10388 11340 11116 11396
rect 11172 11340 11182 11396
rect 11452 11284 11508 11452
rect 12562 11340 12572 11396
rect 12628 11340 16716 11396
rect 16772 11340 18844 11396
rect 18900 11340 18910 11396
rect 22418 11340 22428 11396
rect 22484 11340 22988 11396
rect 23044 11340 23054 11396
rect 24210 11340 24220 11396
rect 24276 11340 26124 11396
rect 26180 11340 26190 11396
rect 28354 11340 28364 11396
rect 28420 11340 31836 11396
rect 31892 11340 31902 11396
rect 37986 11340 37996 11396
rect 38052 11340 46956 11396
rect 47012 11340 47022 11396
rect 47618 11340 47628 11396
rect 47684 11340 49308 11396
rect 49364 11340 49374 11396
rect 52210 11340 52220 11396
rect 52276 11340 54236 11396
rect 54292 11340 54302 11396
rect 10658 11228 10668 11284
rect 10724 11228 11508 11284
rect 11666 11228 11676 11284
rect 11732 11228 14700 11284
rect 14756 11228 14766 11284
rect 17266 11228 17276 11284
rect 17332 11228 18620 11284
rect 18676 11228 18686 11284
rect 25890 11228 25900 11284
rect 25956 11228 27020 11284
rect 27076 11228 27086 11284
rect 27234 11228 27244 11284
rect 27300 11228 28700 11284
rect 28756 11228 28766 11284
rect 30482 11228 30492 11284
rect 30548 11228 30558 11284
rect 30706 11228 30716 11284
rect 30772 11228 31724 11284
rect 31780 11228 35084 11284
rect 35140 11228 35150 11284
rect 9314 11116 9324 11172
rect 9380 11116 17892 11172
rect 18022 11116 18060 11172
rect 18116 11116 18126 11172
rect 9650 11004 9660 11060
rect 9716 11004 14028 11060
rect 14084 11004 14094 11060
rect 14354 11004 14364 11060
rect 14420 11004 15036 11060
rect 15092 11004 15102 11060
rect 6626 10892 6636 10948
rect 6692 10892 6972 10948
rect 7028 10892 7308 10948
rect 7364 10892 8092 10948
rect 8148 10892 11564 10948
rect 11620 10892 11630 10948
rect 13794 10892 13804 10948
rect 13860 10892 14812 10948
rect 14868 10892 17612 10948
rect 17668 10892 17678 10948
rect 17836 10836 17892 11116
rect 30492 11060 30548 11228
rect 31798 11116 31836 11172
rect 31892 11116 31902 11172
rect 35522 11116 35532 11172
rect 35588 11116 36204 11172
rect 36260 11116 36270 11172
rect 37874 11116 37884 11172
rect 37940 11116 38556 11172
rect 38612 11116 38622 11172
rect 23874 11004 23884 11060
rect 23940 11004 30548 11060
rect 42802 11004 42812 11060
rect 42868 11004 43428 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 43372 10948 43428 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 18610 10892 18620 10948
rect 18676 10892 19068 10948
rect 19124 10892 19134 10948
rect 20738 10892 20748 10948
rect 20804 10892 29148 10948
rect 29204 10892 29214 10948
rect 29362 10892 29372 10948
rect 29428 10892 31388 10948
rect 31444 10892 31454 10948
rect 31602 10892 31612 10948
rect 31668 10892 31706 10948
rect 43362 10892 43372 10948
rect 43428 10892 43438 10948
rect 20748 10836 20804 10892
rect 7074 10780 7084 10836
rect 7140 10780 8540 10836
rect 8596 10780 8606 10836
rect 10098 10780 10108 10836
rect 10164 10780 17556 10836
rect 17714 10780 17724 10836
rect 17780 10780 20524 10836
rect 20580 10780 20804 10836
rect 24098 10780 24108 10836
rect 24164 10780 24332 10836
rect 24388 10780 24398 10836
rect 24546 10780 24556 10836
rect 24612 10780 27580 10836
rect 27636 10780 27646 10836
rect 28354 10780 28364 10836
rect 28420 10780 35644 10836
rect 35700 10780 35710 10836
rect 39890 10780 39900 10836
rect 39956 10780 41356 10836
rect 41412 10780 41692 10836
rect 41748 10780 41758 10836
rect 17500 10724 17556 10780
rect 10658 10668 10668 10724
rect 10724 10668 11676 10724
rect 11732 10668 12908 10724
rect 12964 10668 12974 10724
rect 14018 10668 14028 10724
rect 14084 10668 17276 10724
rect 17332 10668 17342 10724
rect 17500 10668 19180 10724
rect 19236 10668 25004 10724
rect 25060 10668 25070 10724
rect 25554 10668 25564 10724
rect 25620 10668 30324 10724
rect 31042 10668 31052 10724
rect 31108 10668 31612 10724
rect 31668 10668 33292 10724
rect 33348 10668 33358 10724
rect 34514 10668 34524 10724
rect 34580 10668 37100 10724
rect 37156 10668 37660 10724
rect 37716 10668 38332 10724
rect 38388 10668 38398 10724
rect 46722 10668 46732 10724
rect 46788 10668 47964 10724
rect 48020 10668 48030 10724
rect 30268 10612 30324 10668
rect 6514 10556 6524 10612
rect 6580 10556 7756 10612
rect 7812 10556 7822 10612
rect 7970 10556 7980 10612
rect 8036 10556 12124 10612
rect 12180 10556 13244 10612
rect 13300 10556 13310 10612
rect 14802 10556 14812 10612
rect 14868 10556 14924 10612
rect 14980 10556 14990 10612
rect 17938 10556 17948 10612
rect 18004 10556 19292 10612
rect 19348 10556 19358 10612
rect 20402 10556 20412 10612
rect 20468 10556 22204 10612
rect 22260 10556 22270 10612
rect 22530 10556 22540 10612
rect 22596 10556 23884 10612
rect 23940 10556 23950 10612
rect 24882 10556 24892 10612
rect 24948 10556 26684 10612
rect 26740 10556 29372 10612
rect 29428 10556 29438 10612
rect 30258 10556 30268 10612
rect 30324 10556 35756 10612
rect 35812 10556 35822 10612
rect 41458 10556 41468 10612
rect 41524 10556 42028 10612
rect 42084 10556 43260 10612
rect 43316 10556 44940 10612
rect 44996 10556 45006 10612
rect 47282 10556 47292 10612
rect 47348 10556 48076 10612
rect 48132 10556 48142 10612
rect 48626 10556 48636 10612
rect 48692 10556 49644 10612
rect 49700 10556 49710 10612
rect 50418 10556 50428 10612
rect 50484 10556 51100 10612
rect 51156 10556 51166 10612
rect 49644 10500 49700 10556
rect 8306 10444 8316 10500
rect 8372 10444 11452 10500
rect 11508 10444 11518 10500
rect 11778 10444 11788 10500
rect 11844 10444 15820 10500
rect 15876 10444 16828 10500
rect 16884 10444 16894 10500
rect 18050 10444 18060 10500
rect 18116 10444 20188 10500
rect 20244 10444 20254 10500
rect 24658 10444 24668 10500
rect 24724 10444 25564 10500
rect 25620 10444 25630 10500
rect 28130 10444 28140 10500
rect 28196 10444 28924 10500
rect 28980 10444 28990 10500
rect 30818 10444 30828 10500
rect 30884 10444 32284 10500
rect 32340 10444 32620 10500
rect 32676 10444 32686 10500
rect 42242 10444 42252 10500
rect 42308 10444 42812 10500
rect 42868 10444 45164 10500
rect 45220 10444 45230 10500
rect 49644 10444 50764 10500
rect 50820 10444 50830 10500
rect 13906 10332 13916 10388
rect 13972 10332 14588 10388
rect 14644 10332 15260 10388
rect 15316 10332 15326 10388
rect 18396 10332 19516 10388
rect 19572 10332 19740 10388
rect 19796 10332 24780 10388
rect 24836 10332 26236 10388
rect 26292 10332 26302 10388
rect 45042 10332 45052 10388
rect 45108 10332 45836 10388
rect 45892 10332 45902 10388
rect 50082 10332 50092 10388
rect 50148 10332 50540 10388
rect 50596 10332 51212 10388
rect 51268 10332 51278 10388
rect 18396 10276 18452 10332
rect 12562 10220 12572 10276
rect 12628 10220 14252 10276
rect 14308 10220 14318 10276
rect 14802 10220 14812 10276
rect 14868 10220 14924 10276
rect 14980 10220 14990 10276
rect 18386 10220 18396 10276
rect 18452 10220 18462 10276
rect 18610 10220 18620 10276
rect 18676 10220 19068 10276
rect 19124 10220 21308 10276
rect 21364 10220 24668 10276
rect 24724 10220 24734 10276
rect 29810 10220 29820 10276
rect 29876 10220 32508 10276
rect 32564 10220 32574 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 12450 10108 12460 10164
rect 12516 10108 13356 10164
rect 13412 10108 13422 10164
rect 14130 10108 14140 10164
rect 14196 10108 14812 10164
rect 14868 10108 14878 10164
rect 16258 10108 16268 10164
rect 16324 10108 23324 10164
rect 23380 10108 24444 10164
rect 24500 10108 24510 10164
rect 6066 9996 6076 10052
rect 6132 9996 9436 10052
rect 9492 9996 11452 10052
rect 11508 9996 11518 10052
rect 14354 9996 14364 10052
rect 14420 9996 15372 10052
rect 15428 9996 15438 10052
rect 16118 9996 16156 10052
rect 16212 9996 16222 10052
rect 20514 9996 20524 10052
rect 20580 9996 23548 10052
rect 23604 9996 23614 10052
rect 24658 9996 24668 10052
rect 24724 9996 27244 10052
rect 27300 9996 27916 10052
rect 27972 9996 27982 10052
rect 33394 9996 33404 10052
rect 33460 9996 39564 10052
rect 39620 9996 41020 10052
rect 41076 9996 41804 10052
rect 41860 9996 41870 10052
rect 43474 9996 43484 10052
rect 43540 9996 44604 10052
rect 44660 9996 44670 10052
rect 5954 9884 5964 9940
rect 6020 9884 9884 9940
rect 9940 9884 11396 9940
rect 13682 9884 13692 9940
rect 13748 9884 20860 9940
rect 20916 9884 20926 9940
rect 22754 9884 22764 9940
rect 22820 9884 23100 9940
rect 23156 9884 25452 9940
rect 25508 9884 25518 9940
rect 26898 9884 26908 9940
rect 26964 9884 27356 9940
rect 27412 9884 27422 9940
rect 31490 9884 31500 9940
rect 31556 9884 31836 9940
rect 31892 9884 31902 9940
rect 35858 9884 35868 9940
rect 35924 9884 37100 9940
rect 37156 9884 37166 9940
rect 38546 9884 38556 9940
rect 38612 9884 38892 9940
rect 38948 9884 38958 9940
rect 11340 9828 11396 9884
rect 27356 9828 27412 9884
rect 7746 9772 7756 9828
rect 7812 9772 8876 9828
rect 8932 9772 10556 9828
rect 10612 9772 10622 9828
rect 11330 9772 11340 9828
rect 11396 9772 12236 9828
rect 12292 9772 12302 9828
rect 12898 9772 12908 9828
rect 12964 9772 14476 9828
rect 14532 9772 14542 9828
rect 15362 9772 15372 9828
rect 15428 9772 17388 9828
rect 17444 9772 17454 9828
rect 21074 9772 21084 9828
rect 21140 9772 21756 9828
rect 21812 9772 21822 9828
rect 24210 9772 24220 9828
rect 24276 9772 25116 9828
rect 25172 9772 25182 9828
rect 26852 9772 27020 9828
rect 27076 9772 27086 9828
rect 27356 9772 28252 9828
rect 28308 9772 28318 9828
rect 28690 9772 28700 9828
rect 28756 9772 34300 9828
rect 34356 9772 35084 9828
rect 35140 9772 35150 9828
rect 37986 9772 37996 9828
rect 38052 9772 46620 9828
rect 46676 9772 46686 9828
rect 26852 9716 26908 9772
rect 9874 9660 9884 9716
rect 9940 9660 12684 9716
rect 12740 9660 13580 9716
rect 13636 9660 13646 9716
rect 14578 9660 14588 9716
rect 14644 9660 15484 9716
rect 15540 9660 15550 9716
rect 18162 9660 18172 9716
rect 18228 9660 18620 9716
rect 18676 9660 18686 9716
rect 22978 9660 22988 9716
rect 23044 9660 26908 9716
rect 33394 9660 33404 9716
rect 33460 9660 39340 9716
rect 39396 9660 40572 9716
rect 40628 9660 40638 9716
rect 50194 9660 50204 9716
rect 50260 9660 51660 9716
rect 51716 9660 51726 9716
rect 3266 9548 3276 9604
rect 3332 9548 11004 9604
rect 11060 9548 11070 9604
rect 12338 9548 12348 9604
rect 12404 9548 13132 9604
rect 13188 9548 13198 9604
rect 13356 9548 16044 9604
rect 16100 9548 25340 9604
rect 25396 9548 25406 9604
rect 32946 9548 32956 9604
rect 33012 9548 36204 9604
rect 36260 9548 36270 9604
rect 42914 9548 42924 9604
rect 42980 9548 43484 9604
rect 43540 9548 43550 9604
rect 13356 9492 13412 9548
rect 6850 9436 6860 9492
rect 6916 9436 6926 9492
rect 9090 9436 9100 9492
rect 9156 9436 13412 9492
rect 15250 9436 15260 9492
rect 15316 9436 16156 9492
rect 16212 9436 16222 9492
rect 17154 9436 17164 9492
rect 17220 9436 18396 9492
rect 18452 9436 18462 9492
rect 21186 9436 21196 9492
rect 21252 9436 24108 9492
rect 24164 9436 24174 9492
rect 6860 9380 6916 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 6860 9324 13692 9380
rect 13748 9324 15036 9380
rect 15092 9324 19684 9380
rect 19628 9268 19684 9324
rect 21196 9268 21252 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 6178 9212 6188 9268
rect 6244 9212 6860 9268
rect 6916 9212 7756 9268
rect 7812 9212 9436 9268
rect 9492 9212 9502 9268
rect 11218 9212 11228 9268
rect 11284 9212 16492 9268
rect 16548 9212 16558 9268
rect 19628 9212 21252 9268
rect 22194 9212 22204 9268
rect 22260 9212 22764 9268
rect 22820 9212 22830 9268
rect 27682 9212 27692 9268
rect 27748 9212 28812 9268
rect 28868 9212 28878 9268
rect 45266 9212 45276 9268
rect 45332 9212 45612 9268
rect 45668 9212 46284 9268
rect 46340 9212 46350 9268
rect 11228 9156 11284 9212
rect 8306 9100 8316 9156
rect 8372 9100 11284 9156
rect 12786 9100 12796 9156
rect 12852 9100 14140 9156
rect 14196 9100 14206 9156
rect 15092 9100 17164 9156
rect 17220 9100 17230 9156
rect 17826 9100 17836 9156
rect 17892 9100 19068 9156
rect 19124 9100 19134 9156
rect 22082 9100 22092 9156
rect 22148 9100 23324 9156
rect 23380 9100 24220 9156
rect 24276 9100 24286 9156
rect 26674 9100 26684 9156
rect 26740 9100 28028 9156
rect 28084 9100 29148 9156
rect 29204 9100 29214 9156
rect 30716 9100 32396 9156
rect 32452 9100 33180 9156
rect 33236 9100 33246 9156
rect 37090 9100 37100 9156
rect 37156 9100 38108 9156
rect 38164 9100 38780 9156
rect 38836 9100 38846 9156
rect 40674 9100 40684 9156
rect 40740 9100 40750 9156
rect 42018 9100 42028 9156
rect 42084 9100 42812 9156
rect 42868 9100 42878 9156
rect 47842 9100 47852 9156
rect 47908 9100 48860 9156
rect 48916 9100 48926 9156
rect 11890 8988 11900 9044
rect 11956 8988 12572 9044
rect 12628 8988 12638 9044
rect 13682 8988 13692 9044
rect 13748 8988 14364 9044
rect 14420 8988 14430 9044
rect 14886 8988 14924 9044
rect 14980 8988 14990 9044
rect 15092 8932 15148 9100
rect 30716 9044 30772 9100
rect 40684 9044 40740 9100
rect 15922 8988 15932 9044
rect 15988 8988 15998 9044
rect 16146 8988 16156 9044
rect 16212 8988 21532 9044
rect 21588 8988 23660 9044
rect 23716 8988 23884 9044
rect 23940 8988 23950 9044
rect 27122 8988 27132 9044
rect 27188 8988 30772 9044
rect 30930 8988 30940 9044
rect 30996 8988 33068 9044
rect 33124 8988 33134 9044
rect 39330 8988 39340 9044
rect 39396 8988 40740 9044
rect 51986 8988 51996 9044
rect 52052 8988 52668 9044
rect 52724 8988 52734 9044
rect 13346 8876 13356 8932
rect 13412 8876 15148 8932
rect 0 8820 800 8848
rect 15932 8820 15988 8988
rect 16482 8876 16492 8932
rect 16548 8876 21868 8932
rect 21924 8876 21934 8932
rect 22082 8876 22092 8932
rect 22148 8876 25228 8932
rect 25284 8876 25294 8932
rect 25666 8876 25676 8932
rect 25732 8876 26460 8932
rect 26516 8876 31836 8932
rect 31892 8876 31902 8932
rect 34626 8876 34636 8932
rect 34692 8876 36204 8932
rect 36260 8876 36270 8932
rect 44594 8876 44604 8932
rect 44660 8876 44940 8932
rect 44996 8876 45006 8932
rect 51538 8876 51548 8932
rect 51604 8876 52556 8932
rect 52612 8876 52622 8932
rect 59200 8820 60000 8848
rect 0 8764 1708 8820
rect 1764 8764 1774 8820
rect 10546 8764 10556 8820
rect 10612 8764 15484 8820
rect 15540 8764 15988 8820
rect 16706 8764 16716 8820
rect 16772 8764 18060 8820
rect 18116 8764 18126 8820
rect 19506 8764 19516 8820
rect 19572 8764 22204 8820
rect 22260 8764 22270 8820
rect 22754 8764 22764 8820
rect 22820 8764 23436 8820
rect 23492 8764 23502 8820
rect 25442 8764 25452 8820
rect 25508 8764 32956 8820
rect 33012 8764 33022 8820
rect 41234 8764 41244 8820
rect 41300 8764 43932 8820
rect 43988 8764 43998 8820
rect 59052 8764 60000 8820
rect 0 8736 800 8764
rect 25452 8708 25508 8764
rect 8642 8652 8652 8708
rect 8708 8652 11004 8708
rect 11060 8652 11070 8708
rect 12338 8652 12348 8708
rect 12404 8652 18172 8708
rect 18228 8652 18238 8708
rect 20514 8652 20524 8708
rect 20580 8652 23660 8708
rect 23716 8652 25508 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 9762 8540 9772 8596
rect 9828 8540 14364 8596
rect 14420 8540 14430 8596
rect 15362 8540 15372 8596
rect 15428 8540 20412 8596
rect 20468 8540 20478 8596
rect 25330 8540 25340 8596
rect 25396 8540 26236 8596
rect 26292 8540 33740 8596
rect 33796 8540 34636 8596
rect 34692 8540 34702 8596
rect 59052 8484 59108 8764
rect 59200 8736 60000 8764
rect 6402 8428 6412 8484
rect 6468 8428 7420 8484
rect 7476 8428 9884 8484
rect 9940 8428 9950 8484
rect 11676 8428 12908 8484
rect 12964 8428 12974 8484
rect 13570 8428 13580 8484
rect 13636 8428 21084 8484
rect 21140 8428 21150 8484
rect 21942 8428 21980 8484
rect 22036 8428 22046 8484
rect 26898 8428 26908 8484
rect 26964 8428 29708 8484
rect 29764 8428 29774 8484
rect 31826 8428 31836 8484
rect 31892 8428 33852 8484
rect 33908 8428 33918 8484
rect 43698 8428 43708 8484
rect 43764 8428 45276 8484
rect 45332 8428 45342 8484
rect 59052 8428 59332 8484
rect 11676 8372 11732 8428
rect 59276 8372 59332 8428
rect 6290 8316 6300 8372
rect 6356 8316 7644 8372
rect 7700 8316 7980 8372
rect 8036 8316 8046 8372
rect 9090 8316 9100 8372
rect 9156 8316 11732 8372
rect 14438 8316 14476 8372
rect 14532 8316 14542 8372
rect 14690 8316 14700 8372
rect 14756 8316 16380 8372
rect 16436 8316 16446 8372
rect 17490 8316 17500 8372
rect 17556 8316 24556 8372
rect 24612 8316 24622 8372
rect 25218 8316 25228 8372
rect 25284 8316 26124 8372
rect 26180 8316 26190 8372
rect 28354 8316 28364 8372
rect 28420 8316 30044 8372
rect 30100 8316 30110 8372
rect 30594 8316 30604 8372
rect 30660 8316 30670 8372
rect 35634 8316 35644 8372
rect 35700 8316 36204 8372
rect 36260 8316 36988 8372
rect 37044 8316 37884 8372
rect 37940 8316 37950 8372
rect 45490 8316 45500 8372
rect 45556 8316 47740 8372
rect 47796 8316 49308 8372
rect 49364 8316 49532 8372
rect 49588 8316 49598 8372
rect 57922 8316 57932 8372
rect 57988 8316 59332 8372
rect 30604 8260 30660 8316
rect 6514 8204 6524 8260
rect 6580 8204 8428 8260
rect 8484 8204 9772 8260
rect 9828 8204 9838 8260
rect 11218 8204 11228 8260
rect 11284 8204 12236 8260
rect 12292 8204 13580 8260
rect 13636 8204 13646 8260
rect 16454 8204 16492 8260
rect 16548 8204 16558 8260
rect 17938 8204 17948 8260
rect 18004 8204 18508 8260
rect 18564 8204 18574 8260
rect 18834 8204 18844 8260
rect 18900 8204 19292 8260
rect 19348 8204 19358 8260
rect 21410 8204 21420 8260
rect 21476 8204 22316 8260
rect 22372 8204 23100 8260
rect 23156 8204 23166 8260
rect 24322 8204 24332 8260
rect 24388 8204 25788 8260
rect 25844 8204 25854 8260
rect 27990 8204 28028 8260
rect 28084 8204 28094 8260
rect 29334 8204 29372 8260
rect 29428 8204 29438 8260
rect 29922 8204 29932 8260
rect 29988 8204 30660 8260
rect 39890 8204 39900 8260
rect 39956 8204 40572 8260
rect 40628 8204 40638 8260
rect 54002 8204 54012 8260
rect 54068 8204 55580 8260
rect 55636 8204 55646 8260
rect 12786 8092 12796 8148
rect 12852 8092 14140 8148
rect 14196 8092 14206 8148
rect 14588 8092 15988 8148
rect 16818 8092 16828 8148
rect 16884 8092 20188 8148
rect 20244 8092 20254 8148
rect 21074 8092 21084 8148
rect 21140 8092 21644 8148
rect 21700 8092 25228 8148
rect 25284 8092 25294 8148
rect 26338 8092 26348 8148
rect 26404 8092 29036 8148
rect 29092 8092 30604 8148
rect 30660 8092 30670 8148
rect 36306 8092 36316 8148
rect 36372 8092 37212 8148
rect 37268 8092 38444 8148
rect 38500 8092 38510 8148
rect 14588 8036 14644 8092
rect 13794 7980 13804 8036
rect 13860 7980 14644 8036
rect 15932 8036 15988 8092
rect 15932 7980 17836 8036
rect 17892 7980 19516 8036
rect 19572 7980 19582 8036
rect 22530 7980 22540 8036
rect 22596 7980 23436 8036
rect 23492 7980 27020 8036
rect 27076 7980 27086 8036
rect 30342 7980 30380 8036
rect 30436 7980 30446 8036
rect 30930 7980 30940 8036
rect 30996 7980 31612 8036
rect 31668 7980 31678 8036
rect 32498 7980 32508 8036
rect 32564 7980 34972 8036
rect 35028 7980 35038 8036
rect 48402 7980 48412 8036
rect 48468 7980 48972 8036
rect 49028 7980 49038 8036
rect 7298 7868 7308 7924
rect 7364 7868 9884 7924
rect 9940 7868 11788 7924
rect 11844 7868 11854 7924
rect 14812 7868 16044 7924
rect 16100 7868 16110 7924
rect 19030 7868 19068 7924
rect 19124 7868 19134 7924
rect 20290 7868 20300 7924
rect 20356 7868 28028 7924
rect 28084 7868 28094 7924
rect 13346 7756 13356 7812
rect 13412 7756 14588 7812
rect 14644 7756 14654 7812
rect 14812 7700 14868 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 15092 7756 17276 7812
rect 17332 7756 17342 7812
rect 27682 7756 27692 7812
rect 27748 7756 31052 7812
rect 31108 7756 31118 7812
rect 11302 7644 11340 7700
rect 11396 7644 11406 7700
rect 13234 7644 13244 7700
rect 13300 7644 14868 7700
rect 15026 7644 15036 7700
rect 15092 7644 15148 7756
rect 16930 7644 16940 7700
rect 16996 7644 25620 7700
rect 25778 7644 25788 7700
rect 25844 7644 27916 7700
rect 27972 7644 27982 7700
rect 28130 7644 28140 7700
rect 28196 7644 30716 7700
rect 30772 7644 30782 7700
rect 36642 7644 36652 7700
rect 36708 7644 37548 7700
rect 37604 7644 37614 7700
rect 25564 7588 25620 7644
rect 13122 7532 13132 7588
rect 13188 7532 13916 7588
rect 13972 7532 13982 7588
rect 14466 7532 14476 7588
rect 14532 7532 15708 7588
rect 15764 7532 15774 7588
rect 16034 7532 16044 7588
rect 16100 7532 20524 7588
rect 20580 7532 20590 7588
rect 24098 7532 24108 7588
rect 24164 7532 25340 7588
rect 25396 7532 25406 7588
rect 25564 7532 28028 7588
rect 28084 7532 28588 7588
rect 28644 7532 28654 7588
rect 30146 7532 30156 7588
rect 30212 7532 36540 7588
rect 36596 7532 36606 7588
rect 13010 7420 13020 7476
rect 13076 7420 13468 7476
rect 13524 7420 15036 7476
rect 15092 7420 15102 7476
rect 15474 7420 15484 7476
rect 15540 7420 16380 7476
rect 16436 7420 16446 7476
rect 20290 7420 20300 7476
rect 20356 7420 20636 7476
rect 20692 7420 24444 7476
rect 24500 7420 24510 7476
rect 27906 7420 27916 7476
rect 27972 7420 28140 7476
rect 28196 7420 28206 7476
rect 29138 7420 29148 7476
rect 29204 7420 30380 7476
rect 30436 7420 30446 7476
rect 30706 7420 30716 7476
rect 30772 7420 32844 7476
rect 32900 7420 32910 7476
rect 33730 7420 33740 7476
rect 33796 7420 34748 7476
rect 34804 7420 34814 7476
rect 38658 7420 38668 7476
rect 38724 7420 39116 7476
rect 39172 7420 39182 7476
rect 44258 7420 44268 7476
rect 44324 7420 45500 7476
rect 45556 7420 46284 7476
rect 46340 7420 46350 7476
rect 49298 7420 49308 7476
rect 49364 7420 51436 7476
rect 51492 7420 51502 7476
rect 10770 7308 10780 7364
rect 10836 7308 15148 7364
rect 16818 7308 16828 7364
rect 16884 7308 17836 7364
rect 17892 7308 18508 7364
rect 18564 7308 24220 7364
rect 24276 7308 24286 7364
rect 34178 7308 34188 7364
rect 34244 7308 34972 7364
rect 35028 7308 35038 7364
rect 35634 7308 35644 7364
rect 35700 7308 37100 7364
rect 37156 7308 37166 7364
rect 37986 7308 37996 7364
rect 38052 7308 43932 7364
rect 43988 7308 45276 7364
rect 45332 7308 45342 7364
rect 7634 7196 7644 7252
rect 7700 7196 10332 7252
rect 10388 7196 13692 7252
rect 13748 7196 13758 7252
rect 15092 7140 15148 7308
rect 16034 7196 16044 7252
rect 16100 7196 18732 7252
rect 18788 7196 18798 7252
rect 19170 7196 19180 7252
rect 19236 7196 21084 7252
rect 21140 7196 21150 7252
rect 25330 7196 25340 7252
rect 25396 7196 28140 7252
rect 28196 7196 28206 7252
rect 28466 7196 28476 7252
rect 28532 7196 30604 7252
rect 30660 7196 30670 7252
rect 37538 7196 37548 7252
rect 37604 7196 38332 7252
rect 38388 7196 38398 7252
rect 41906 7196 41916 7252
rect 41972 7196 42476 7252
rect 42532 7196 42542 7252
rect 46162 7196 46172 7252
rect 46228 7196 47964 7252
rect 48020 7196 49196 7252
rect 49252 7196 49262 7252
rect 11442 7084 11452 7140
rect 11508 7084 14924 7140
rect 14980 7084 14990 7140
rect 15092 7084 16492 7140
rect 16548 7084 16940 7140
rect 16996 7084 17006 7140
rect 18946 7084 18956 7140
rect 19012 7084 27916 7140
rect 27972 7084 27982 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 7746 6972 7756 7028
rect 7812 6972 10948 7028
rect 11666 6972 11676 7028
rect 11732 6972 19180 7028
rect 19236 6972 19246 7028
rect 20178 6972 20188 7028
rect 20244 6972 21308 7028
rect 21364 6972 23436 7028
rect 23492 6972 24276 7028
rect 26562 6972 26572 7028
rect 26628 6972 27356 7028
rect 27412 6972 27422 7028
rect 10892 6916 10948 6972
rect 6738 6860 6748 6916
rect 6804 6860 8204 6916
rect 8260 6860 8270 6916
rect 10892 6860 11732 6916
rect 12898 6860 12908 6916
rect 12964 6860 15148 6916
rect 15204 6860 15214 6916
rect 16370 6860 16380 6916
rect 16436 6860 17500 6916
rect 17556 6860 17566 6916
rect 19394 6860 19404 6916
rect 19460 6860 19852 6916
rect 19908 6860 19918 6916
rect 11676 6804 11732 6860
rect 24220 6804 24276 6972
rect 24434 6860 24444 6916
rect 24500 6860 27692 6916
rect 27748 6860 27758 6916
rect 33170 6860 33180 6916
rect 33236 6860 35196 6916
rect 35252 6860 35262 6916
rect 7298 6748 7308 6804
rect 7364 6748 7980 6804
rect 8036 6748 9548 6804
rect 9604 6748 9614 6804
rect 10444 6748 11452 6804
rect 11508 6748 11518 6804
rect 11666 6748 11676 6804
rect 11732 6748 13244 6804
rect 13300 6748 13310 6804
rect 15092 6748 21196 6804
rect 21252 6748 21262 6804
rect 22502 6748 22540 6804
rect 22596 6748 22606 6804
rect 24220 6748 26684 6804
rect 26740 6748 26750 6804
rect 27234 6748 27244 6804
rect 27300 6748 33516 6804
rect 33572 6748 33582 6804
rect 40226 6748 40236 6804
rect 40292 6748 41188 6804
rect 49858 6748 49868 6804
rect 49924 6748 50540 6804
rect 50596 6748 50606 6804
rect 10444 6692 10500 6748
rect 15092 6692 15148 6748
rect 41132 6692 41188 6748
rect 8988 6636 10500 6692
rect 10658 6636 10668 6692
rect 10724 6636 11116 6692
rect 11172 6636 14028 6692
rect 14084 6636 15148 6692
rect 16566 6636 16604 6692
rect 16660 6636 16670 6692
rect 18386 6636 18396 6692
rect 18452 6636 19964 6692
rect 20020 6636 21308 6692
rect 21364 6636 21980 6692
rect 22036 6636 22046 6692
rect 26684 6636 32284 6692
rect 32340 6636 32350 6692
rect 37986 6636 37996 6692
rect 38052 6636 40908 6692
rect 40964 6636 40974 6692
rect 41132 6636 41356 6692
rect 41412 6636 43484 6692
rect 43540 6636 43550 6692
rect 50372 6636 50652 6692
rect 50708 6636 50718 6692
rect 8988 6468 9044 6636
rect 9874 6524 9884 6580
rect 9940 6524 12684 6580
rect 12740 6524 12750 6580
rect 13346 6524 13356 6580
rect 13412 6524 13692 6580
rect 13748 6524 13758 6580
rect 16258 6524 16268 6580
rect 16324 6524 18284 6580
rect 18340 6524 24108 6580
rect 24164 6524 24174 6580
rect 26684 6468 26740 6636
rect 27794 6524 27804 6580
rect 27860 6524 28812 6580
rect 28868 6524 28878 6580
rect 32162 6524 32172 6580
rect 32228 6524 34076 6580
rect 34132 6524 34142 6580
rect 36530 6524 36540 6580
rect 36596 6524 38444 6580
rect 38500 6524 38510 6580
rect 41906 6524 41916 6580
rect 41972 6524 46732 6580
rect 46788 6524 46798 6580
rect 8978 6412 8988 6468
rect 9044 6412 9054 6468
rect 9650 6412 9660 6468
rect 9716 6412 12908 6468
rect 12964 6412 12974 6468
rect 15250 6412 15260 6468
rect 15316 6412 15932 6468
rect 15988 6412 15998 6468
rect 16370 6412 16380 6468
rect 16436 6412 19068 6468
rect 19124 6412 19134 6468
rect 19628 6412 21420 6468
rect 21476 6412 21486 6468
rect 26674 6412 26684 6468
rect 26740 6412 26750 6468
rect 26898 6412 26908 6468
rect 26964 6412 27244 6468
rect 27300 6412 27468 6468
rect 27524 6412 27534 6468
rect 31490 6412 31500 6468
rect 31556 6412 33852 6468
rect 33908 6412 33918 6468
rect 34514 6412 34524 6468
rect 34580 6412 40348 6468
rect 40404 6412 40414 6468
rect 11330 6300 11340 6356
rect 11396 6300 18956 6356
rect 19012 6300 19022 6356
rect 19628 6244 19684 6412
rect 50372 6356 50428 6636
rect 47954 6300 47964 6356
rect 48020 6300 50428 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 7746 6188 7756 6244
rect 7812 6188 11788 6244
rect 11844 6188 12628 6244
rect 15362 6188 15372 6244
rect 15428 6188 16156 6244
rect 16212 6188 16222 6244
rect 16818 6188 16828 6244
rect 16884 6188 19684 6244
rect 21410 6188 21420 6244
rect 21476 6188 21756 6244
rect 21812 6188 21822 6244
rect 23426 6188 23436 6244
rect 23492 6188 35644 6244
rect 35700 6188 36316 6244
rect 36372 6188 37324 6244
rect 37380 6188 37390 6244
rect 12572 6132 12628 6188
rect 9762 6076 9772 6132
rect 9828 6076 12124 6132
rect 12180 6076 12190 6132
rect 12534 6076 12572 6132
rect 12628 6076 12638 6132
rect 16034 6076 16044 6132
rect 16100 6076 18396 6132
rect 18452 6076 18462 6132
rect 19366 6076 19404 6132
rect 19460 6076 19470 6132
rect 24546 6076 24556 6132
rect 24612 6076 26796 6132
rect 26852 6076 34076 6132
rect 34132 6076 34142 6132
rect 9426 5964 9436 6020
rect 9492 5964 15036 6020
rect 15092 5964 15102 6020
rect 15586 5964 15596 6020
rect 15652 5964 16380 6020
rect 16436 5964 16446 6020
rect 16818 5964 16828 6020
rect 16884 5964 16894 6020
rect 17266 5964 17276 6020
rect 17332 5964 18060 6020
rect 18116 5964 18126 6020
rect 19170 5964 19180 6020
rect 19236 5964 22092 6020
rect 22148 5964 22158 6020
rect 22978 5964 22988 6020
rect 23044 5964 25228 6020
rect 25284 5964 25294 6020
rect 25778 5964 25788 6020
rect 25844 5964 27020 6020
rect 27076 5964 27580 6020
rect 27636 5964 27646 6020
rect 29698 5964 29708 6020
rect 29764 5964 30604 6020
rect 30660 5964 30670 6020
rect 32162 5964 32172 6020
rect 32228 5964 32620 6020
rect 32676 5964 32686 6020
rect 35186 5964 35196 6020
rect 35252 5964 42140 6020
rect 42196 5964 42206 6020
rect 46498 5964 46508 6020
rect 46564 5964 47180 6020
rect 47236 5964 47246 6020
rect 16828 5908 16884 5964
rect 7186 5852 7196 5908
rect 7252 5852 10220 5908
rect 10276 5852 10286 5908
rect 12114 5852 12124 5908
rect 12180 5852 17500 5908
rect 17556 5852 17566 5908
rect 20626 5852 20636 5908
rect 20692 5852 23100 5908
rect 23156 5852 23166 5908
rect 27346 5852 27356 5908
rect 27412 5852 27804 5908
rect 27860 5852 29148 5908
rect 29204 5852 29214 5908
rect 31154 5852 31164 5908
rect 31220 5852 31948 5908
rect 32004 5852 32014 5908
rect 33628 5852 33964 5908
rect 34020 5852 34030 5908
rect 33628 5796 33684 5852
rect 10098 5740 10108 5796
rect 10164 5740 13692 5796
rect 13748 5740 13758 5796
rect 14438 5740 14476 5796
rect 14532 5740 14542 5796
rect 15810 5740 15820 5796
rect 15876 5740 19068 5796
rect 19124 5740 21532 5796
rect 21588 5740 21598 5796
rect 26450 5740 26460 5796
rect 26516 5740 28476 5796
rect 28532 5740 28542 5796
rect 31714 5740 31724 5796
rect 31780 5740 33628 5796
rect 33684 5740 33694 5796
rect 13794 5628 13804 5684
rect 13860 5628 18396 5684
rect 18452 5628 18462 5684
rect 18834 5628 18844 5684
rect 18900 5628 20860 5684
rect 20916 5628 20926 5684
rect 22082 5628 22092 5684
rect 22148 5628 26012 5684
rect 26068 5628 26078 5684
rect 27682 5628 27692 5684
rect 27748 5628 31836 5684
rect 31892 5628 31902 5684
rect 36082 5628 36092 5684
rect 36148 5628 38892 5684
rect 38948 5628 39452 5684
rect 39508 5628 39518 5684
rect 10658 5516 10668 5572
rect 10724 5516 13916 5572
rect 13972 5516 13982 5572
rect 15138 5516 15148 5572
rect 15204 5516 18620 5572
rect 18676 5516 18686 5572
rect 19030 5516 19068 5572
rect 19124 5516 19134 5572
rect 20402 5516 20412 5572
rect 20468 5516 24332 5572
rect 24388 5516 24398 5572
rect 26226 5516 26236 5572
rect 26292 5516 28252 5572
rect 28308 5516 29036 5572
rect 29092 5516 32340 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 13916 5460 13972 5516
rect 13916 5404 17948 5460
rect 18004 5404 18014 5460
rect 21298 5404 21308 5460
rect 21364 5404 31276 5460
rect 31332 5404 31342 5460
rect 32284 5348 32340 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 59200 5460 60000 5488
rect 58146 5404 58156 5460
rect 58212 5404 60000 5460
rect 59200 5376 60000 5404
rect 12674 5292 12684 5348
rect 12740 5292 13468 5348
rect 13524 5292 13534 5348
rect 14242 5292 14252 5348
rect 14308 5292 14318 5348
rect 16482 5292 16492 5348
rect 16548 5292 16940 5348
rect 16996 5292 17006 5348
rect 19618 5292 19628 5348
rect 19684 5292 23324 5348
rect 23380 5292 26348 5348
rect 26404 5292 26414 5348
rect 29922 5292 29932 5348
rect 29988 5292 31500 5348
rect 31556 5292 32060 5348
rect 32116 5292 32126 5348
rect 32284 5292 35420 5348
rect 35476 5292 35486 5348
rect 9202 5180 9212 5236
rect 9268 5180 11564 5236
rect 11620 5180 11630 5236
rect 13234 5180 13244 5236
rect 13300 5180 13692 5236
rect 13748 5180 13758 5236
rect 14252 5124 14308 5292
rect 14466 5180 14476 5236
rect 14532 5180 14924 5236
rect 14980 5180 14990 5236
rect 15138 5180 15148 5236
rect 15204 5180 16716 5236
rect 16772 5180 16782 5236
rect 21186 5180 21196 5236
rect 21252 5180 22540 5236
rect 22596 5180 24332 5236
rect 24388 5180 24398 5236
rect 26562 5180 26572 5236
rect 26628 5180 27356 5236
rect 27412 5180 27422 5236
rect 31602 5180 31612 5236
rect 31668 5180 33292 5236
rect 33348 5180 33358 5236
rect 41122 5180 41132 5236
rect 41188 5180 42812 5236
rect 42868 5180 45388 5236
rect 45444 5180 46172 5236
rect 46228 5180 46238 5236
rect 8530 5068 8540 5124
rect 8596 5068 12236 5124
rect 12292 5068 13580 5124
rect 13636 5068 13646 5124
rect 14252 5068 18116 5124
rect 18274 5068 18284 5124
rect 18340 5068 21308 5124
rect 21364 5068 21374 5124
rect 29026 5068 29036 5124
rect 29092 5068 29708 5124
rect 29764 5068 29774 5124
rect 32386 5068 32396 5124
rect 32452 5068 33740 5124
rect 33796 5068 33806 5124
rect 39778 5068 39788 5124
rect 39844 5068 40684 5124
rect 40740 5068 40750 5124
rect 42578 5068 42588 5124
rect 42644 5068 43372 5124
rect 43428 5068 45164 5124
rect 45220 5068 46396 5124
rect 46452 5068 46462 5124
rect 18060 5012 18116 5068
rect 11778 4956 11788 5012
rect 11844 4956 16604 5012
rect 16660 4956 16670 5012
rect 18060 4956 24444 5012
rect 24500 4956 26572 5012
rect 26628 4956 26638 5012
rect 29250 4956 29260 5012
rect 29316 4956 30044 5012
rect 30100 4956 32172 5012
rect 32228 4956 32238 5012
rect 33068 4956 33180 5012
rect 33236 4956 33246 5012
rect 39666 4956 39676 5012
rect 39732 4956 41244 5012
rect 41300 4956 41310 5012
rect 33068 4900 33124 4956
rect 12562 4844 12572 4900
rect 12628 4844 14140 4900
rect 14196 4844 18060 4900
rect 18116 4844 19292 4900
rect 19348 4844 19358 4900
rect 20962 4844 20972 4900
rect 21028 4844 26124 4900
rect 26180 4844 26190 4900
rect 26338 4844 26348 4900
rect 26404 4844 27356 4900
rect 27412 4844 27422 4900
rect 28364 4844 33124 4900
rect 28364 4788 28420 4844
rect 59200 4788 60000 4816
rect 13346 4732 13356 4788
rect 13412 4732 13916 4788
rect 13972 4732 13982 4788
rect 14466 4732 14476 4788
rect 14532 4732 15876 4788
rect 18274 4732 18284 4788
rect 18340 4732 19516 4788
rect 19572 4732 19582 4788
rect 20850 4732 20860 4788
rect 20916 4732 28420 4788
rect 28578 4732 28588 4788
rect 28644 4732 28924 4788
rect 28980 4732 30940 4788
rect 30996 4732 33180 4788
rect 33236 4732 33246 4788
rect 58146 4732 58156 4788
rect 58212 4732 60000 4788
rect 15820 4676 15876 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 59200 4704 60000 4732
rect 12674 4620 12684 4676
rect 12740 4620 15596 4676
rect 15652 4620 15662 4676
rect 15820 4620 19180 4676
rect 19236 4620 19246 4676
rect 24210 4620 24220 4676
rect 24276 4620 26516 4676
rect 26460 4564 26516 4620
rect 10098 4508 10108 4564
rect 10164 4508 10668 4564
rect 10724 4508 10734 4564
rect 10882 4508 10892 4564
rect 10948 4508 11788 4564
rect 11844 4508 13692 4564
rect 13748 4508 13758 4564
rect 16034 4508 16044 4564
rect 16100 4508 16380 4564
rect 16436 4508 16446 4564
rect 16594 4508 16604 4564
rect 16660 4508 17724 4564
rect 17780 4508 17790 4564
rect 18498 4508 18508 4564
rect 18564 4508 26236 4564
rect 26292 4508 26302 4564
rect 26460 4508 27244 4564
rect 27300 4508 27310 4564
rect 27458 4508 27468 4564
rect 27524 4508 34524 4564
rect 34580 4508 34590 4564
rect 10434 4396 10444 4452
rect 10500 4396 11900 4452
rect 11956 4396 11966 4452
rect 14130 4396 14140 4452
rect 14196 4396 15260 4452
rect 15316 4396 21420 4452
rect 21476 4396 21486 4452
rect 12226 4284 12236 4340
rect 12292 4284 12908 4340
rect 12964 4284 14812 4340
rect 14868 4284 16268 4340
rect 16324 4284 17164 4340
rect 17220 4284 17230 4340
rect 19282 4284 19292 4340
rect 19348 4284 19964 4340
rect 20020 4284 20030 4340
rect 23986 4284 23996 4340
rect 24052 4284 26684 4340
rect 26740 4284 29148 4340
rect 29204 4284 29214 4340
rect 40338 4284 40348 4340
rect 40404 4284 41132 4340
rect 41188 4284 41198 4340
rect 15474 4172 15484 4228
rect 15540 4172 18956 4228
rect 19012 4172 19022 4228
rect 19170 4172 19180 4228
rect 19236 4172 21756 4228
rect 21812 4172 21822 4228
rect 25554 4172 25564 4228
rect 25620 4172 28700 4228
rect 28756 4172 29484 4228
rect 29540 4172 29550 4228
rect 30146 4172 30156 4228
rect 30212 4172 32172 4228
rect 32228 4172 32238 4228
rect 59200 4116 60000 4144
rect 14690 4060 14700 4116
rect 14756 4060 22428 4116
rect 22484 4060 23436 4116
rect 23492 4060 23502 4116
rect 58146 4060 58156 4116
rect 58212 4060 60000 4116
rect 59200 4032 60000 4060
rect 14242 3948 14252 4004
rect 14308 3948 19180 4004
rect 19236 3948 19246 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 13346 3836 13356 3892
rect 13412 3836 14476 3892
rect 14532 3836 14542 3892
rect 16482 3836 16492 3892
rect 16548 3836 20972 3892
rect 21028 3836 21038 3892
rect 21410 3836 21420 3892
rect 21476 3836 29708 3892
rect 29764 3836 30828 3892
rect 30884 3836 33180 3892
rect 33236 3836 33246 3892
rect 17042 3724 17052 3780
rect 17108 3724 20300 3780
rect 20356 3724 20366 3780
rect 11554 3612 11564 3668
rect 11620 3612 14140 3668
rect 14196 3612 14206 3668
rect 15092 3556 15148 3668
rect 15204 3612 15214 3668
rect 16006 3612 16044 3668
rect 16100 3612 16110 3668
rect 17714 3612 17724 3668
rect 17780 3612 18396 3668
rect 18452 3612 18462 3668
rect 18946 3612 18956 3668
rect 19012 3612 22764 3668
rect 22820 3612 22830 3668
rect 27346 3612 27356 3668
rect 27412 3612 34076 3668
rect 34132 3612 34142 3668
rect 51762 3612 51772 3668
rect 51828 3612 52892 3668
rect 52948 3612 52958 3668
rect 13458 3500 13468 3556
rect 13524 3500 15148 3556
rect 15586 3500 15596 3556
rect 15652 3500 16716 3556
rect 16772 3500 16782 3556
rect 19170 3500 19180 3556
rect 19236 3500 23548 3556
rect 23604 3500 23614 3556
rect 27794 3500 27804 3556
rect 27860 3500 28476 3556
rect 28532 3500 31612 3556
rect 31668 3500 31678 3556
rect 59200 3444 60000 3472
rect 10658 3388 10668 3444
rect 10724 3388 14252 3444
rect 14308 3388 14588 3444
rect 14644 3388 14654 3444
rect 19842 3388 19852 3444
rect 19908 3388 23212 3444
rect 23268 3388 23278 3444
rect 29474 3388 29484 3444
rect 29540 3388 32396 3444
rect 32452 3388 32462 3444
rect 43698 3388 43708 3444
rect 43764 3388 44940 3444
rect 44996 3388 45006 3444
rect 58380 3388 60000 3444
rect 58380 3332 58436 3388
rect 59200 3360 60000 3388
rect 7746 3276 7756 3332
rect 7812 3276 8428 3332
rect 10770 3276 10780 3332
rect 10836 3276 19068 3332
rect 19124 3276 19134 3332
rect 19292 3276 22036 3332
rect 22978 3276 22988 3332
rect 23044 3276 32732 3332
rect 32788 3276 32798 3332
rect 58146 3276 58156 3332
rect 58212 3276 58436 3332
rect 8372 2996 8428 3276
rect 19292 3220 19348 3276
rect 8978 3164 8988 3220
rect 9044 3164 15820 3220
rect 15876 3164 15886 3220
rect 17826 3164 17836 3220
rect 17892 3164 19348 3220
rect 21980 3220 22036 3276
rect 21980 3164 39116 3220
rect 39172 3164 39182 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 11666 3052 11676 3108
rect 11732 3052 17276 3108
rect 17332 3052 17342 3108
rect 20402 3052 20412 3108
rect 20468 3052 38780 3108
rect 38836 3052 38846 3108
rect 8372 2940 15932 2996
rect 15988 2940 19516 2996
rect 19572 2940 19582 2996
rect 8306 2828 8316 2884
rect 8372 2772 8428 2884
rect 15362 2828 15372 2884
rect 15428 2828 29484 2884
rect 29540 2828 29550 2884
rect 59200 2772 60000 2800
rect 8372 2716 14924 2772
rect 14980 2716 14990 2772
rect 15138 2716 15148 2772
rect 15204 2716 18956 2772
rect 19012 2716 19022 2772
rect 57698 2716 57708 2772
rect 57764 2716 60000 2772
rect 59200 2688 60000 2716
rect 17714 2604 17724 2660
rect 17780 2604 36876 2660
rect 36932 2604 36942 2660
rect 11330 2492 11340 2548
rect 11396 2492 18060 2548
rect 18116 2492 18126 2548
rect 16930 2380 16940 2436
rect 16996 2380 32508 2436
rect 32564 2380 32574 2436
rect 23492 2268 24668 2324
rect 24724 2268 24734 2324
rect 23492 2212 23548 2268
rect 14914 2156 14924 2212
rect 14980 2156 23548 2212
rect 18834 1596 18844 1652
rect 18900 1596 26908 1652
rect 26964 1596 26974 1652
rect 18050 1484 18060 1540
rect 18116 1484 39004 1540
rect 39060 1484 39070 1540
rect 7858 1372 7868 1428
rect 7924 1372 30380 1428
rect 30436 1372 30446 1428
<< via3 >>
rect 28140 57148 28196 57204
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 30380 56028 30436 56084
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 15820 55580 15876 55636
rect 28588 55580 28644 55636
rect 20972 55468 21028 55524
rect 28700 55468 28756 55524
rect 27468 55020 27524 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19516 53788 19572 53844
rect 22316 53788 22372 53844
rect 20748 53452 20804 53508
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 19404 53228 19460 53284
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 21196 52444 21252 52500
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19628 51772 19684 51828
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 23660 51436 23716 51492
rect 18396 51324 18452 51380
rect 22988 51212 23044 51268
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 16604 50876 16660 50932
rect 20972 50764 21028 50820
rect 18956 50652 19012 50708
rect 22316 50540 22372 50596
rect 25564 50540 25620 50596
rect 43036 50540 43092 50596
rect 28476 50428 28532 50484
rect 30492 50316 30548 50372
rect 19516 50204 19572 50260
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 18956 50092 19012 50148
rect 18620 49980 18676 50036
rect 23996 49868 24052 49924
rect 21196 49532 21252 49588
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 21756 49084 21812 49140
rect 16604 48972 16660 49028
rect 23212 48748 23268 48804
rect 31388 48748 31444 48804
rect 43036 48748 43092 48804
rect 27356 48636 27412 48692
rect 30492 48636 30548 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 22764 48524 22820 48580
rect 23324 48524 23380 48580
rect 22876 48412 22932 48468
rect 22652 48188 22708 48244
rect 18508 48076 18564 48132
rect 25564 48076 25620 48132
rect 20748 47964 20804 48020
rect 23996 47852 24052 47908
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 22876 47740 22932 47796
rect 22988 47628 23044 47684
rect 22764 47516 22820 47572
rect 18396 47180 18452 47236
rect 18620 47180 18676 47236
rect 23492 47180 23548 47236
rect 27356 47180 27412 47236
rect 18508 47068 18564 47124
rect 19068 47068 19124 47124
rect 19404 47068 19460 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 13580 46956 13636 47012
rect 19292 46956 19348 47012
rect 23548 46956 23604 47012
rect 22652 46844 22708 46900
rect 23884 46732 23940 46788
rect 19068 46620 19124 46676
rect 30828 46620 30884 46676
rect 23212 46508 23268 46564
rect 20748 46396 20804 46452
rect 26796 46396 26852 46452
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 21980 46172 22036 46228
rect 27804 46172 27860 46228
rect 28028 46172 28084 46228
rect 15932 45836 15988 45892
rect 19068 45612 19124 45668
rect 28028 45612 28084 45668
rect 26908 45500 26964 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 19516 45276 19572 45332
rect 17052 45164 17108 45220
rect 28588 45052 28644 45108
rect 34412 45052 34468 45108
rect 16044 44940 16100 44996
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 17052 44604 17108 44660
rect 15820 44492 15876 44548
rect 19292 44492 19348 44548
rect 13580 44268 13636 44324
rect 18060 44044 18116 44100
rect 18844 43932 18900 43988
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 18732 43708 18788 43764
rect 15708 43484 15764 43540
rect 26348 43484 26404 43540
rect 28140 43260 28196 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 15932 43036 15988 43092
rect 27580 43036 27636 43092
rect 28476 43036 28532 43092
rect 34300 43036 34356 43092
rect 27020 42924 27076 42980
rect 18844 42700 18900 42756
rect 19628 42700 19684 42756
rect 28140 42588 28196 42644
rect 31612 42476 31668 42532
rect 27020 42364 27076 42420
rect 27804 42364 27860 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 19628 42252 19684 42308
rect 26796 42252 26852 42308
rect 27580 42252 27636 42308
rect 34300 42252 34356 42308
rect 15260 42140 15316 42196
rect 23548 42140 23604 42196
rect 14252 42028 14308 42084
rect 26572 42028 26628 42084
rect 28700 41804 28756 41860
rect 15260 41580 15316 41636
rect 16044 41580 16100 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19404 41356 19460 41412
rect 26572 41356 26628 41412
rect 27020 41244 27076 41300
rect 25228 41132 25284 41188
rect 27804 41132 27860 41188
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 20748 40684 20804 40740
rect 18956 40572 19012 40628
rect 18732 40460 18788 40516
rect 19516 40348 19572 40404
rect 19292 40124 19348 40180
rect 19516 40124 19572 40180
rect 18956 40012 19012 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 23436 39788 23492 39844
rect 25228 39788 25284 39844
rect 20188 39676 20244 39732
rect 23884 39676 23940 39732
rect 30828 39564 30884 39620
rect 25116 39340 25172 39396
rect 31612 39340 31668 39396
rect 19068 39228 19124 39284
rect 20860 39228 20916 39284
rect 21756 39228 21812 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 20860 38668 20916 38724
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 26348 38332 26404 38388
rect 15932 38220 15988 38276
rect 34412 38108 34468 38164
rect 19628 37996 19684 38052
rect 19404 37772 19460 37828
rect 25116 37660 25172 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 18620 37548 18676 37604
rect 21980 37548 22036 37604
rect 14252 37324 14308 37380
rect 30268 37100 30324 37156
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 27468 36876 27524 36932
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 18620 36540 18676 36596
rect 20188 36428 20244 36484
rect 19292 36204 19348 36260
rect 15708 36092 15764 36148
rect 19628 36092 19684 36148
rect 20188 36092 20244 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 25116 35980 25172 36036
rect 18060 35308 18116 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 31388 35084 31444 35140
rect 19404 34748 19460 34804
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 30380 33292 30436 33348
rect 19404 32844 19460 32900
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 30380 32732 30436 32788
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 23996 31836 24052 31892
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 30268 31276 30324 31332
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 43596 27132 43652 27188
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 43596 26236 43652 26292
rect 29036 26124 29092 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 29036 25676 29092 25732
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 16156 23772 16212 23828
rect 22204 23772 22260 23828
rect 21980 23548 22036 23604
rect 22204 23548 22260 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 14924 23436 14980 23492
rect 26124 22988 26180 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19516 22652 19572 22708
rect 26908 22428 26964 22484
rect 12908 22092 12964 22148
rect 30716 21980 30772 22036
rect 46284 21980 46340 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 22428 21868 22484 21924
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 20524 21532 20580 21588
rect 24556 21308 24612 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 20524 20972 20580 21028
rect 13692 20860 13748 20916
rect 22428 20748 22484 20804
rect 28028 20524 28084 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 28588 20188 28644 20244
rect 34412 20188 34468 20244
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 32956 19180 33012 19236
rect 7980 19068 8036 19124
rect 11340 18844 11396 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 16716 18620 16772 18676
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 14476 18396 14532 18452
rect 21980 18396 22036 18452
rect 27580 18396 27636 18452
rect 7980 18172 8036 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 20636 17836 20692 17892
rect 24556 17836 24612 17892
rect 30716 17836 30772 17892
rect 27244 17612 27300 17668
rect 14252 17388 14308 17444
rect 14588 17388 14644 17444
rect 27356 17388 27412 17444
rect 27916 17388 27972 17444
rect 10108 17276 10164 17332
rect 20188 17276 20244 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 27244 17052 27300 17108
rect 8316 16828 8372 16884
rect 34412 16716 34468 16772
rect 29372 16604 29428 16660
rect 34860 16604 34916 16660
rect 17164 16492 17220 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 18172 16380 18228 16436
rect 20188 16380 20244 16436
rect 32956 16380 33012 16436
rect 33516 16380 33572 16436
rect 15372 16268 15428 16324
rect 27580 16268 27636 16324
rect 31836 16044 31892 16100
rect 16604 15820 16660 15876
rect 27356 15820 27412 15876
rect 15372 15708 15428 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 24332 15260 24388 15316
rect 28700 15260 28756 15316
rect 15036 15148 15092 15204
rect 12908 14924 12964 14980
rect 16044 14924 16100 14980
rect 28700 14924 28756 14980
rect 33516 14924 33572 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 46508 14812 46564 14868
rect 23436 14476 23492 14532
rect 46508 14252 46564 14308
rect 19628 14140 19684 14196
rect 27916 14140 27972 14196
rect 46284 14140 46340 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 17164 14028 17220 14084
rect 23548 13916 23604 13972
rect 18172 13580 18228 13636
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 14252 13020 14308 13076
rect 14476 13020 14532 13076
rect 26124 12908 26180 12964
rect 10108 12796 10164 12852
rect 27916 12684 27972 12740
rect 20524 12572 20580 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 13580 12460 13636 12516
rect 19628 12236 19684 12292
rect 28588 12236 28644 12292
rect 7980 12124 8036 12180
rect 20636 11788 20692 11844
rect 34860 11788 34916 11844
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 11452 11676 11508 11732
rect 18172 11676 18228 11732
rect 28364 11676 28420 11732
rect 10668 11564 10724 11620
rect 11228 11564 11284 11620
rect 10780 11452 10836 11508
rect 19068 11452 19124 11508
rect 43484 11452 43540 11508
rect 16716 11340 16772 11396
rect 28364 11340 28420 11396
rect 31836 11340 31892 11396
rect 17276 11228 17332 11284
rect 18060 11116 18116 11172
rect 14364 11004 14420 11060
rect 31836 11116 31892 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 29372 10892 29428 10948
rect 31612 10892 31668 10948
rect 24332 10780 24388 10836
rect 10668 10668 10724 10724
rect 17276 10668 17332 10724
rect 14812 10556 14868 10612
rect 22540 10556 22596 10612
rect 8316 10444 8372 10500
rect 11452 10444 11508 10500
rect 19516 10332 19572 10388
rect 12572 10220 12628 10276
rect 14812 10220 14868 10276
rect 18396 10220 18452 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 23324 10108 23380 10164
rect 16156 9996 16212 10052
rect 23548 9996 23604 10052
rect 26908 9884 26964 9940
rect 31836 9884 31892 9940
rect 43484 9548 43540 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 15036 9324 15092 9380
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 14364 8988 14420 9044
rect 14924 8988 14980 9044
rect 18172 8652 18228 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 14364 8540 14420 8596
rect 21980 8428 22036 8484
rect 14476 8316 14532 8372
rect 26124 8316 26180 8372
rect 16492 8204 16548 8260
rect 28028 8204 28084 8260
rect 29372 8204 29428 8260
rect 30380 7980 30436 8036
rect 31612 7980 31668 8036
rect 19068 7868 19124 7924
rect 14588 7756 14644 7812
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 11340 7644 11396 7700
rect 15036 7644 15092 7700
rect 14476 7532 14532 7588
rect 16044 7532 16100 7588
rect 14924 7084 14980 7140
rect 16940 7084 16996 7140
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 23436 6972 23492 7028
rect 16380 6860 16436 6916
rect 19404 6860 19460 6916
rect 22540 6748 22596 6804
rect 16604 6636 16660 6692
rect 21980 6636 22036 6692
rect 19068 6412 19124 6468
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 11788 6188 11844 6244
rect 16828 6188 16884 6244
rect 12572 6076 12628 6132
rect 18396 6076 18452 6132
rect 19404 6076 19460 6132
rect 14476 5740 14532 5796
rect 19068 5516 19124 5572
rect 29036 5516 29092 5572
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 23324 5292 23380 5348
rect 16604 4956 16660 5012
rect 14476 4732 14532 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 19180 4620 19236 4676
rect 11788 4508 11844 4564
rect 16380 4508 16436 4564
rect 19180 4172 19236 4228
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 14476 3836 14532 3892
rect 16044 3612 16100 3668
rect 16716 3500 16772 3556
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 16940 2380 16996 2436
rect 18060 1484 18116 1540
rect 30380 1372 30436 1428
<< metal4 >>
rect 28140 57204 28196 57214
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 15820 55636 15876 55646
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 13580 47012 13636 47022
rect 13580 44324 13636 46956
rect 15820 44548 15876 55580
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19516 53844 19572 53854
rect 19404 53284 19460 53294
rect 18396 51380 18452 51390
rect 16604 50932 16660 50942
rect 16604 49028 16660 50876
rect 16604 48962 16660 48972
rect 18396 47236 18452 51324
rect 18956 50708 19012 50718
rect 18956 50148 19012 50652
rect 18956 50082 19012 50092
rect 18620 50036 18676 50046
rect 18396 47170 18452 47180
rect 18508 48132 18564 48142
rect 18508 47124 18564 48076
rect 18620 47236 18676 49980
rect 18620 47170 18676 47180
rect 18508 47058 18564 47068
rect 19068 47124 19124 47134
rect 19068 46676 19124 47068
rect 19404 47124 19460 53228
rect 19516 50260 19572 53788
rect 19808 53340 20128 54852
rect 20972 55524 21028 55534
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19516 50194 19572 50204
rect 19628 51828 19684 51838
rect 19404 47058 19460 47068
rect 19068 46610 19124 46620
rect 19292 47012 19348 47022
rect 15820 44482 15876 44492
rect 15932 45892 15988 45902
rect 13580 44258 13636 44268
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 15708 43540 15764 43550
rect 15260 42196 15316 42206
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 14252 42084 14308 42094
rect 14252 37380 14308 42028
rect 15260 41636 15316 42140
rect 15260 41570 15316 41580
rect 14252 37314 14308 37324
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 15708 36148 15764 43484
rect 15932 43092 15988 45836
rect 19068 45668 19124 45678
rect 17052 45220 17108 45230
rect 15932 38276 15988 43036
rect 16044 44996 16100 45006
rect 16044 41636 16100 44940
rect 17052 44660 17108 45164
rect 17052 44594 17108 44604
rect 16044 41570 16100 41580
rect 18060 44100 18116 44110
rect 15932 38210 15988 38220
rect 15708 36082 15764 36092
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 18060 35364 18116 44044
rect 18844 43988 18900 43998
rect 18732 43764 18788 43774
rect 18732 40516 18788 43708
rect 18844 42756 18900 43932
rect 18844 42690 18900 42700
rect 18732 40450 18788 40460
rect 18956 40628 19012 40638
rect 18956 40068 19012 40572
rect 18956 40002 19012 40012
rect 19068 39284 19124 45612
rect 19068 39218 19124 39228
rect 19292 44548 19348 46956
rect 19292 40180 19348 44492
rect 19516 45332 19572 45342
rect 18620 37604 18676 37614
rect 18620 36596 18676 37548
rect 18620 36530 18676 36540
rect 19292 36260 19348 40124
rect 19404 41412 19460 41422
rect 19404 37828 19460 41356
rect 19516 40404 19572 45276
rect 19628 42756 19684 51772
rect 19628 42690 19684 42700
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 20748 53508 20804 53518
rect 20748 48020 20804 53452
rect 20972 50820 21028 55468
rect 27468 55076 27524 55086
rect 22316 53844 22372 53854
rect 20972 50754 21028 50764
rect 21196 52500 21252 52510
rect 21196 49588 21252 52444
rect 22316 50596 22372 53788
rect 23660 51492 23716 51502
rect 22316 50530 22372 50540
rect 22988 51268 23044 51278
rect 21196 49522 21252 49532
rect 20748 47954 20804 47964
rect 21756 49140 21812 49150
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19516 40180 19572 40348
rect 19516 40114 19572 40124
rect 19628 42308 19684 42318
rect 19404 37762 19460 37772
rect 19628 38052 19684 42252
rect 19292 36194 19348 36204
rect 19628 36148 19684 37996
rect 19628 36082 19684 36092
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 20748 46452 20804 46462
rect 20748 40740 20804 46396
rect 20748 40674 20804 40684
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 18060 35298 18116 35308
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 20188 39732 20244 39742
rect 20188 36484 20244 39676
rect 20860 39284 20916 39294
rect 20860 38724 20916 39228
rect 21756 39284 21812 49084
rect 22764 48580 22820 48590
rect 22652 48244 22708 48254
rect 22652 46900 22708 48188
rect 22764 47572 22820 48524
rect 22876 48468 22932 48478
rect 22876 47796 22932 48412
rect 22876 47730 22932 47740
rect 22988 47684 23044 51212
rect 23212 48804 23268 48814
rect 23212 48538 23268 48748
rect 22988 47618 23044 47628
rect 23100 48482 23268 48538
rect 23324 48580 23380 48590
rect 22764 47506 22820 47516
rect 23100 47278 23156 48482
rect 23324 47278 23380 48524
rect 23100 47222 23268 47278
rect 23324 47236 23548 47278
rect 23324 47222 23492 47236
rect 22652 46834 22708 46844
rect 23212 46564 23268 47222
rect 23492 47170 23548 47180
rect 23660 47098 23716 51436
rect 25564 50596 25620 50606
rect 23548 47042 23716 47098
rect 23996 49924 24052 49934
rect 23996 47908 24052 49868
rect 25564 48132 25620 50540
rect 25564 48066 25620 48076
rect 27356 48692 27412 48702
rect 23548 47012 23604 47042
rect 23548 46946 23604 46956
rect 23212 46498 23268 46508
rect 23884 46788 23940 46798
rect 21756 39218 21812 39228
rect 21980 46228 22036 46238
rect 20860 38658 20916 38668
rect 21980 37604 22036 46172
rect 23548 42196 23604 42206
rect 23548 40438 23604 42140
rect 23436 40382 23604 40438
rect 23436 39844 23492 40382
rect 23436 39778 23492 39788
rect 23884 39732 23940 46732
rect 23884 39666 23940 39676
rect 21980 37538 22036 37548
rect 20188 36148 20244 36428
rect 20188 36082 20244 36092
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19404 34804 19460 34814
rect 19404 32900 19460 34748
rect 19404 32834 19460 32844
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 19808 31388 20128 32900
rect 23996 31892 24052 47852
rect 27356 47236 27412 48636
rect 27356 47170 27412 47180
rect 26796 46452 26852 46462
rect 26348 43540 26404 43550
rect 25228 41188 25284 41198
rect 25228 39844 25284 41132
rect 25228 39778 25284 39788
rect 25116 39396 25172 39406
rect 25116 37716 25172 39340
rect 26348 38388 26404 43484
rect 26796 42308 26852 46396
rect 26908 45556 26964 45566
rect 26964 45500 27076 45556
rect 26908 45490 26964 45500
rect 27020 42980 27076 45500
rect 27020 42914 27076 42924
rect 26796 42242 26852 42252
rect 27020 42420 27076 42430
rect 26572 42084 26628 42094
rect 26572 41412 26628 42028
rect 26572 41346 26628 41356
rect 27020 41300 27076 42364
rect 27020 41234 27076 41244
rect 26348 38322 26404 38332
rect 25116 36036 25172 37660
rect 27468 36932 27524 55020
rect 27804 46228 27860 46238
rect 27580 43092 27636 43102
rect 27580 42308 27636 43036
rect 27580 42242 27636 42252
rect 27804 42420 27860 46172
rect 28028 46228 28084 46238
rect 28028 45668 28084 46172
rect 28028 45602 28084 45612
rect 28140 43316 28196 57148
rect 30380 56084 30436 56094
rect 28588 55636 28644 55646
rect 28140 42644 28196 43260
rect 28476 50484 28532 50494
rect 28476 43092 28532 50428
rect 28588 45108 28644 55580
rect 28588 45042 28644 45052
rect 28700 55524 28756 55534
rect 28476 43026 28532 43036
rect 28140 42578 28196 42588
rect 27804 41188 27860 42364
rect 28700 41860 28756 55468
rect 28700 41794 28756 41804
rect 27804 41122 27860 41132
rect 27468 36866 27524 36876
rect 30268 37156 30324 37166
rect 25116 35970 25172 35980
rect 23996 31826 24052 31836
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 30268 31332 30324 37100
rect 30380 33348 30436 56028
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 30492 50372 30548 50382
rect 30492 48692 30548 50316
rect 35168 49420 35488 50932
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 30492 48626 30548 48636
rect 31388 48804 31444 48814
rect 30828 46676 30884 46686
rect 30828 39620 30884 46620
rect 30828 39554 30884 39564
rect 31388 35140 31444 48748
rect 35168 47852 35488 49364
rect 43036 50596 43092 50606
rect 43036 48804 43092 50540
rect 43036 48738 43092 48748
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 34412 45108 34468 45118
rect 34300 43092 34356 43102
rect 31612 42532 31668 42542
rect 31612 39396 31668 42476
rect 34300 42308 34356 43036
rect 34300 42242 34356 42252
rect 31612 39330 31668 39340
rect 34412 38164 34468 45052
rect 34412 38098 34468 38108
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 31388 35074 31444 35084
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 30380 32788 30436 33292
rect 30380 32722 30436 32732
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 30268 31266 30324 31276
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 16156 23828 16212 23838
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 14924 23492 14980 23502
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 12908 22148 12964 22158
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 7980 19124 8036 19134
rect 7980 18228 8036 19068
rect 7980 12180 8036 18172
rect 11340 18900 11396 18910
rect 10108 17332 10164 17342
rect 7980 12114 8036 12124
rect 8316 16884 8372 16894
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 8316 10500 8372 16828
rect 10108 12852 10164 17276
rect 10108 12786 10164 12796
rect 10668 11620 10724 11630
rect 10668 10724 10724 11564
rect 10780 11620 11284 11638
rect 10780 11582 11228 11620
rect 10780 11508 10836 11582
rect 11228 11554 11284 11564
rect 10780 11442 10836 11452
rect 10668 10658 10724 10668
rect 8316 10434 8372 10444
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 11340 7700 11396 18844
rect 12908 14980 12964 22092
rect 13692 20916 13748 20926
rect 13692 15148 13748 20860
rect 14476 18452 14532 18462
rect 12908 14914 12964 14924
rect 13580 15092 13748 15148
rect 14252 17444 14308 17454
rect 13580 12516 13636 15092
rect 14252 13076 14308 17388
rect 14252 13010 14308 13020
rect 14476 13076 14532 18396
rect 14476 13010 14532 13020
rect 14588 17444 14644 17454
rect 13580 12450 13636 12460
rect 11452 11732 11508 11742
rect 11452 10500 11508 11676
rect 11452 10434 11508 10444
rect 14364 11060 14420 11070
rect 11340 7634 11396 7644
rect 12572 10276 12628 10286
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 11788 6244 11844 6254
rect 11788 4564 11844 6188
rect 12572 6132 12628 10220
rect 14364 9044 14420 11004
rect 14364 8596 14420 8988
rect 14364 7318 14420 8540
rect 14476 8372 14532 8382
rect 14476 7588 14532 8316
rect 14588 7812 14644 17388
rect 14812 10612 14868 10622
rect 14812 10276 14868 10556
rect 14812 10210 14868 10220
rect 14924 9044 14980 23436
rect 15372 16324 15428 16334
rect 15372 15764 15428 16268
rect 15372 15698 15428 15708
rect 15036 15204 15092 15214
rect 15036 9380 15092 15148
rect 15036 9314 15092 9324
rect 16044 14980 16100 14990
rect 14924 8978 14980 8988
rect 14588 7746 14644 7756
rect 15036 7700 15092 7710
rect 14476 7522 14532 7532
rect 14924 7644 15036 7678
rect 14924 7622 15092 7644
rect 14364 7262 14532 7318
rect 12572 6066 12628 6076
rect 11788 4498 11844 4508
rect 14476 5796 14532 7262
rect 14924 7140 14980 7622
rect 14924 7074 14980 7084
rect 16044 7588 16100 14924
rect 16156 10052 16212 23772
rect 19808 23548 20128 25060
rect 29036 26180 29092 26190
rect 29036 25732 29092 26124
rect 22204 23828 22260 23838
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19516 22708 19572 22718
rect 16716 18676 16772 18686
rect 16380 18620 16716 18658
rect 16380 18602 16772 18620
rect 16380 15148 16436 18602
rect 17164 16548 17220 16558
rect 16604 15876 16660 15886
rect 16380 15092 16548 15148
rect 16156 9986 16212 9996
rect 16492 8260 16548 15092
rect 16492 8194 16548 8204
rect 14476 4788 14532 5740
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 14476 3892 14532 4732
rect 14476 3826 14532 3836
rect 16044 3668 16100 7532
rect 16380 6916 16436 6926
rect 16380 4564 16436 6860
rect 16604 6692 16660 15820
rect 17164 14084 17220 16492
rect 17164 14018 17220 14028
rect 18172 16436 18228 16446
rect 18172 13636 18228 16380
rect 18172 13570 18228 13580
rect 18172 11732 18228 11742
rect 16604 5012 16660 6636
rect 16604 4946 16660 4956
rect 16716 11396 16772 11406
rect 16716 6238 16772 11340
rect 17276 11284 17332 11294
rect 17276 10724 17332 11228
rect 17276 10658 17332 10668
rect 18060 11172 18116 11182
rect 16940 7140 16996 7150
rect 16828 6244 16884 6254
rect 16716 6188 16828 6238
rect 16716 6182 16884 6188
rect 16380 4498 16436 4508
rect 16044 3602 16100 3612
rect 16716 3556 16772 6182
rect 16828 6178 16884 6182
rect 16716 3490 16772 3500
rect 16940 2436 16996 7084
rect 16940 2370 16996 2380
rect 18060 1540 18116 11116
rect 18172 8708 18228 11676
rect 19068 11508 19124 11518
rect 18172 8642 18228 8652
rect 18396 10276 18452 10286
rect 18396 6132 18452 10220
rect 19068 7924 19124 11452
rect 19516 10388 19572 22652
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 21980 23604 22036 23614
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 20524 21588 20580 21598
rect 20524 21028 20580 21532
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20188 17332 20244 17342
rect 20188 16436 20244 17276
rect 20188 16370 20244 16380
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19628 14196 19684 14206
rect 19628 12292 19684 14140
rect 19628 12226 19684 12236
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 20524 12628 20580 20972
rect 21980 18452 22036 23548
rect 22204 23604 22260 23772
rect 22204 23538 22260 23548
rect 26124 23044 26180 23054
rect 22428 21924 22484 21934
rect 22428 20804 22484 21868
rect 22428 20738 22484 20748
rect 24556 21364 24612 21374
rect 21980 18386 22036 18396
rect 20524 12562 20580 12572
rect 20636 17892 20692 17902
rect 19516 10322 19572 10332
rect 19808 11004 20128 12516
rect 20636 11844 20692 17836
rect 24556 17892 24612 21308
rect 24556 17826 24612 17836
rect 24332 15316 24388 15326
rect 20636 11778 20692 11788
rect 23436 14532 23492 14542
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19068 7858 19124 7868
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 22540 10612 22596 10622
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19404 6916 19460 6926
rect 18396 6066 18452 6076
rect 19068 6468 19124 6478
rect 19068 5572 19124 6412
rect 19404 6132 19460 6860
rect 19404 6066 19460 6076
rect 19808 6300 20128 7812
rect 21980 8484 22036 8494
rect 21980 6692 22036 8428
rect 22540 6804 22596 10556
rect 22540 6738 22596 6748
rect 23324 10164 23380 10174
rect 21980 6626 22036 6636
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19068 5506 19124 5516
rect 19808 4732 20128 6244
rect 23324 5348 23380 10108
rect 23436 7028 23492 14476
rect 23548 13972 23604 13982
rect 23548 10052 23604 13916
rect 24332 10836 24388 15260
rect 24332 10770 24388 10780
rect 26124 12964 26180 22988
rect 23548 9986 23604 9996
rect 26124 8372 26180 12908
rect 26908 22484 26964 22494
rect 26908 9940 26964 22428
rect 28028 20580 28084 20590
rect 27580 18452 27636 18462
rect 27244 17668 27300 17678
rect 27244 17108 27300 17612
rect 27244 17042 27300 17052
rect 27356 17444 27412 17454
rect 27356 15876 27412 17388
rect 27580 16324 27636 18396
rect 27580 16258 27636 16268
rect 27916 17444 27972 17454
rect 27356 15810 27412 15820
rect 27916 14196 27972 17388
rect 27916 12740 27972 14140
rect 27916 12674 27972 12684
rect 26908 9874 26964 9884
rect 26124 8306 26180 8316
rect 28028 8260 28084 20524
rect 28588 20244 28644 20254
rect 28588 12292 28644 20188
rect 28700 15316 28756 15326
rect 28700 14980 28756 15260
rect 28700 14914 28756 14924
rect 28588 12226 28644 12236
rect 28364 11732 28420 11742
rect 28364 11396 28420 11676
rect 28364 11330 28420 11340
rect 28028 8194 28084 8204
rect 23436 6962 23492 6972
rect 29036 5572 29092 25676
rect 35168 25900 35488 27412
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 43596 27188 43652 27198
rect 43596 26292 43652 27132
rect 43596 26226 43652 26236
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 30716 22036 30772 22046
rect 30716 17892 30772 21980
rect 35168 21196 35488 22708
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 34412 20244 34468 20254
rect 30716 17826 30772 17836
rect 32956 19236 33012 19246
rect 29372 16660 29428 16670
rect 29372 10948 29428 16604
rect 32956 16436 33012 19180
rect 34412 16772 34468 20188
rect 34412 16706 34468 16716
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 34860 16660 34916 16670
rect 32956 16370 33012 16380
rect 33516 16436 33572 16446
rect 31836 16100 31892 16110
rect 31836 11396 31892 16044
rect 33516 14980 33572 16380
rect 33516 14914 33572 14924
rect 34860 11844 34916 16604
rect 34860 11778 34916 11788
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 46284 22036 46340 22046
rect 46284 14196 46340 21980
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 46508 14868 46564 14878
rect 46508 14308 46564 14812
rect 46508 14242 46564 14252
rect 46284 14130 46340 14140
rect 50528 14140 50848 15652
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 31836 11172 31892 11340
rect 29372 8260 29428 10892
rect 29372 8194 29428 8204
rect 31612 10948 31668 10958
rect 29036 5506 29092 5516
rect 30380 8036 30436 8046
rect 23324 5282 23380 5292
rect 19180 4676 19236 4686
rect 19180 4228 19236 4620
rect 19180 4162 19236 4172
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 18060 1474 18116 1484
rect 30380 1428 30436 7980
rect 31612 8036 31668 10892
rect 31836 9940 31892 11116
rect 31836 9874 31892 9884
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 31612 7970 31668 7980
rect 35168 8652 35488 10164
rect 43484 11508 43540 11518
rect 43484 9604 43540 11452
rect 43484 9538 43540 9548
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 30380 1362 30436 1372
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1373_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1374_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1375_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1376_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1377_
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1378_
timestamp 1698431365
transform 1 0 10752 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1379_
timestamp 1698431365
transform -1 0 10976 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1380_
timestamp 1698431365
transform -1 0 11984 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1381_
timestamp 1698431365
transform -1 0 22064 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1382_
timestamp 1698431365
transform -1 0 20160 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1383_
timestamp 1698431365
transform 1 0 10528 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1384_
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1385_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1386_
timestamp 1698431365
transform 1 0 23520 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1387_
timestamp 1698431365
transform -1 0 12880 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1388_
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1389_
timestamp 1698431365
transform -1 0 15456 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1390_
timestamp 1698431365
transform 1 0 8960 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1391_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12208 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1392_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1393_
timestamp 1698431365
transform -1 0 30016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1394_
timestamp 1698431365
transform -1 0 29680 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1395_
timestamp 1698431365
transform -1 0 30576 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1396_
timestamp 1698431365
transform 1 0 30912 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1397_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32480 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1398_
timestamp 1698431365
transform -1 0 30912 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1399_
timestamp 1698431365
transform 1 0 12880 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1400_
timestamp 1698431365
transform 1 0 11648 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1401_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1402_
timestamp 1698431365
transform 1 0 17584 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1403_
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1404_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26768 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1405_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1406_
timestamp 1698431365
transform -1 0 29568 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1407_
timestamp 1698431365
transform -1 0 30912 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1408_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30688 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1409_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1410_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32480 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1411_
timestamp 1698431365
transform -1 0 10752 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1412_
timestamp 1698431365
transform -1 0 8960 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1413_
timestamp 1698431365
transform 1 0 8400 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1414_
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1415_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12544 0 1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1416_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29904 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1417_
timestamp 1698431365
transform 1 0 32256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1418_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39872 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1419_
timestamp 1698431365
transform -1 0 8288 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1420_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1421_
timestamp 1698431365
transform 1 0 9520 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1422_
timestamp 1698431365
transform 1 0 6496 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1423_
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1424_
timestamp 1698431365
transform 1 0 9408 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1425_
timestamp 1698431365
transform -1 0 12768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1426_
timestamp 1698431365
transform -1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1427_
timestamp 1698431365
transform 1 0 7504 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1428_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1429_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1430_
timestamp 1698431365
transform -1 0 12544 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1431_
timestamp 1698431365
transform 1 0 5600 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1432_
timestamp 1698431365
transform 1 0 6272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1433_
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1434_
timestamp 1698431365
transform -1 0 10976 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1435_
timestamp 1698431365
transform -1 0 11536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1436_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1437_
timestamp 1698431365
transform -1 0 14784 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1438_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1439_
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1440_
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1441_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1442_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1443_
timestamp 1698431365
transform -1 0 6720 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698431365
transform -1 0 6608 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1445_
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1446_
timestamp 1698431365
transform -1 0 10416 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1447_
timestamp 1698431365
transform 1 0 6160 0 -1 15680
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1448_
timestamp 1698431365
transform 1 0 14784 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1449_
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1450_
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1451_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1452_
timestamp 1698431365
transform -1 0 37744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1453_
timestamp 1698431365
transform 1 0 30800 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1454_
timestamp 1698431365
transform -1 0 35056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1455_
timestamp 1698431365
transform 1 0 35392 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1456_
timestamp 1698431365
transform -1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1457_
timestamp 1698431365
transform -1 0 36400 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1458_
timestamp 1698431365
transform -1 0 35616 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1459_
timestamp 1698431365
transform -1 0 34496 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 34384 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1461_
timestamp 1698431365
transform 1 0 38304 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1462_
timestamp 1698431365
transform 1 0 38752 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1463_
timestamp 1698431365
transform -1 0 32144 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698431365
transform 1 0 38416 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1465_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1466_
timestamp 1698431365
transform -1 0 39984 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1467_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1468_
timestamp 1698431365
transform -1 0 39424 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1469_
timestamp 1698431365
transform 1 0 37072 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1470_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38528 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1471_
timestamp 1698431365
transform -1 0 40096 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1472_
timestamp 1698431365
transform 1 0 36736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1473_
timestamp 1698431365
transform 1 0 37184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1474_
timestamp 1698431365
transform -1 0 40544 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1475_
timestamp 1698431365
transform 1 0 38416 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1476_
timestamp 1698431365
transform 1 0 39312 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1477_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38528 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1478_
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1480_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30800 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698431365
transform -1 0 30352 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1482_
timestamp 1698431365
transform -1 0 39872 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1483_
timestamp 1698431365
transform 1 0 38752 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1698431365
transform 1 0 38752 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1485_
timestamp 1698431365
transform -1 0 45024 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1486_
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1698431365
transform 1 0 11760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1488_
timestamp 1698431365
transform 1 0 12656 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1489_
timestamp 1698431365
transform -1 0 26992 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1490_
timestamp 1698431365
transform -1 0 25984 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1491_
timestamp 1698431365
transform -1 0 7616 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1492_
timestamp 1698431365
transform 1 0 7504 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1493_
timestamp 1698431365
transform -1 0 10976 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1494_
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1495_
timestamp 1698431365
transform 1 0 5488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1496_
timestamp 1698431365
transform 1 0 6720 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1497_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24976 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1498_
timestamp 1698431365
transform 1 0 16128 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1499_
timestamp 1698431365
transform 1 0 27104 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1500_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1501_
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1502_
timestamp 1698431365
transform -1 0 30016 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1503_
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1504_
timestamp 1698431365
transform 1 0 8400 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1505_
timestamp 1698431365
transform 1 0 11424 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1506_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16016 0 1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1507_
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1508_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1509_
timestamp 1698431365
transform 1 0 10080 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1510_
timestamp 1698431365
transform 1 0 25648 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1511_
timestamp 1698431365
transform 1 0 14448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1512_
timestamp 1698431365
transform -1 0 19488 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1513_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32368 0 -1 9408
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1514_
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1515_
timestamp 1698431365
transform 1 0 6944 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1516_
timestamp 1698431365
transform 1 0 6832 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1698431365
transform -1 0 7280 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1518_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1519_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25648 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1520_
timestamp 1698431365
transform -1 0 12096 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1521_
timestamp 1698431365
transform 1 0 10416 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1522_
timestamp 1698431365
transform 1 0 11872 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1523_
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1524_
timestamp 1698431365
transform -1 0 10304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1698431365
transform 1 0 24304 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1526_
timestamp 1698431365
transform -1 0 27776 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1527_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1528_
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1529_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1530_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1531_
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1532_
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1533_
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1534_
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1535_
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1536_
timestamp 1698431365
transform 1 0 29568 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1537_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 1 9408
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1538_
timestamp 1698431365
transform -1 0 42672 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1539_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1540_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6608 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1541_
timestamp 1698431365
transform -1 0 15904 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1542_
timestamp 1698431365
transform -1 0 17024 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1543_
timestamp 1698431365
transform -1 0 7280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1544_
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1545_
timestamp 1698431365
transform -1 0 8288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1546_
timestamp 1698431365
transform 1 0 9968 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1547_
timestamp 1698431365
transform -1 0 12992 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1548_
timestamp 1698431365
transform 1 0 10528 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1549_
timestamp 1698431365
transform 1 0 6048 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1550_
timestamp 1698431365
transform 1 0 12320 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1551_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1552_
timestamp 1698431365
transform -1 0 9184 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1553_
timestamp 1698431365
transform 1 0 10192 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1554_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1555_
timestamp 1698431365
transform 1 0 14000 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1556_
timestamp 1698431365
transform 1 0 7840 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1557_
timestamp 1698431365
transform -1 0 15008 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1558_
timestamp 1698431365
transform 1 0 9184 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1559_
timestamp 1698431365
transform 1 0 12432 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1560_
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1561_
timestamp 1698431365
transform 1 0 13440 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1562_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1563_
timestamp 1698431365
transform -1 0 9520 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1564_
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1565_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17024 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1566_
timestamp 1698431365
transform 1 0 9184 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1567_
timestamp 1698431365
transform -1 0 6944 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1568_
timestamp 1698431365
transform -1 0 8400 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1569_
timestamp 1698431365
transform -1 0 15456 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1570_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1571_
timestamp 1698431365
transform -1 0 15792 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1572_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18928 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1573_
timestamp 1698431365
transform 1 0 43120 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1574_
timestamp 1698431365
transform 1 0 43680 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1575_
timestamp 1698431365
transform 1 0 45808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1576_
timestamp 1698431365
transform -1 0 39872 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1577_
timestamp 1698431365
transform -1 0 40432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1578_
timestamp 1698431365
transform 1 0 12096 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1579_
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1580_
timestamp 1698431365
transform 1 0 10752 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1581_
timestamp 1698431365
transform -1 0 22288 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1582_
timestamp 1698431365
transform -1 0 20832 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1583_
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_4  _1584_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1585_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1586_
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1587_
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1588_
timestamp 1698431365
transform -1 0 16240 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1589_
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1590_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10416 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1591_
timestamp 1698431365
transform 1 0 8400 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1592_
timestamp 1698431365
transform -1 0 11424 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1593_
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1594_
timestamp 1698431365
transform -1 0 15344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1595_
timestamp 1698431365
transform 1 0 13664 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1596_
timestamp 1698431365
transform 1 0 19152 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1597_
timestamp 1698431365
transform -1 0 20496 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1598_
timestamp 1698431365
transform 1 0 19264 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1599_
timestamp 1698431365
transform 1 0 35392 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1600_
timestamp 1698431365
transform 1 0 38640 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1601_
timestamp 1698431365
transform 1 0 39200 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1602_
timestamp 1698431365
transform -1 0 41440 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1603_
timestamp 1698431365
transform 1 0 39312 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1604_
timestamp 1698431365
transform 1 0 39984 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1605_
timestamp 1698431365
transform 1 0 8288 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1606_
timestamp 1698431365
transform 1 0 13552 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1607_
timestamp 1698431365
transform 1 0 21392 0 -1 4704
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1608_
timestamp 1698431365
transform -1 0 27104 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1609_
timestamp 1698431365
transform 1 0 20048 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1611_
timestamp 1698431365
transform 1 0 18928 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1612_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1613_
timestamp 1698431365
transform 1 0 18368 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1614_
timestamp 1698431365
transform 1 0 19152 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1615_
timestamp 1698431365
transform 1 0 17024 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1616_
timestamp 1698431365
transform 1 0 17136 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1617_
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1618_
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1619_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1620_
timestamp 1698431365
transform 1 0 14336 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1621_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1622_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 -1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1623_
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1624_
timestamp 1698431365
transform -1 0 36736 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1625_
timestamp 1698431365
transform -1 0 35952 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1626_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1627_
timestamp 1698431365
transform -1 0 43792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1628_
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform -1 0 20160 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1630_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1631_
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1632_
timestamp 1698431365
transform 1 0 22400 0 1 4704
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1633_
timestamp 1698431365
transform 1 0 18928 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1634_
timestamp 1698431365
transform -1 0 20048 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1635_
timestamp 1698431365
transform 1 0 9968 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1636_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1637_
timestamp 1698431365
transform -1 0 20384 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1638_
timestamp 1698431365
transform -1 0 8400 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1639_
timestamp 1698431365
transform -1 0 8624 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1640_
timestamp 1698431365
transform 1 0 14560 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1641_
timestamp 1698431365
transform 1 0 19152 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1642_
timestamp 1698431365
transform -1 0 22624 0 -1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1643_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22624 0 -1 14112
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1644_
timestamp 1698431365
transform -1 0 39760 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1645_
timestamp 1698431365
transform 1 0 10416 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1646_
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1647_
timestamp 1698431365
transform 1 0 11200 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1648_
timestamp 1698431365
transform -1 0 15344 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1649_
timestamp 1698431365
transform 1 0 12096 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1650_
timestamp 1698431365
transform 1 0 7392 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1651_
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1652_
timestamp 1698431365
transform 1 0 13664 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1653_
timestamp 1698431365
transform 1 0 18032 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1654_
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1655_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1656_
timestamp 1698431365
transform -1 0 13888 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1657_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1658_
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1659_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1660_
timestamp 1698431365
transform 1 0 10752 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1661_
timestamp 1698431365
transform 1 0 9968 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1662_
timestamp 1698431365
transform -1 0 16016 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1663_
timestamp 1698431365
transform -1 0 14448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1664_
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform -1 0 16240 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1666_
timestamp 1698431365
transform -1 0 15008 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1667_
timestamp 1698431365
transform -1 0 15344 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1668_
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1671_
timestamp 1698431365
transform -1 0 15344 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1672_
timestamp 1698431365
transform -1 0 18368 0 1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1673_
timestamp 1698431365
transform 1 0 37856 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1674_
timestamp 1698431365
transform 1 0 41328 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1675_
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1676_
timestamp 1698431365
transform 1 0 42000 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1677_
timestamp 1698431365
transform -1 0 42336 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1678_
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1679_
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1680_
timestamp 1698431365
transform 1 0 10976 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1681_
timestamp 1698431365
transform 1 0 23296 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1682_
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1683_
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1684_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30016 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1685_
timestamp 1698431365
transform -1 0 22736 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1686_
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1687_
timestamp 1698431365
transform 1 0 30016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1688_
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1689_
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1690_
timestamp 1698431365
transform 1 0 25648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1691_
timestamp 1698431365
transform 1 0 30464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1692_
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1693_
timestamp 1698431365
transform -1 0 34384 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1694_
timestamp 1698431365
transform -1 0 34720 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1695_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1696_
timestamp 1698431365
transform 1 0 42672 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1697_
timestamp 1698431365
transform 1 0 41328 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1698_
timestamp 1698431365
transform 1 0 45024 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1699_
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1700_
timestamp 1698431365
transform 1 0 40544 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1701_
timestamp 1698431365
transform 1 0 12096 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1702_
timestamp 1698431365
transform 1 0 17920 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1703_
timestamp 1698431365
transform 1 0 17360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1704_
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1705_
timestamp 1698431365
transform 1 0 17472 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1706_
timestamp 1698431365
transform 1 0 14672 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1707_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1708_
timestamp 1698431365
transform 1 0 14896 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1709_
timestamp 1698431365
transform 1 0 10416 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1710_
timestamp 1698431365
transform 1 0 15456 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1711_
timestamp 1698431365
transform 1 0 16128 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1712_
timestamp 1698431365
transform 1 0 16352 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1713_
timestamp 1698431365
transform 1 0 35952 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1714_
timestamp 1698431365
transform 1 0 38192 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1715_
timestamp 1698431365
transform 1 0 36848 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1716_
timestamp 1698431365
transform 1 0 38416 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1717_
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1718_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10192 0 -1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1719_
timestamp 1698431365
transform 1 0 13440 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1720_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1721_
timestamp 1698431365
transform -1 0 20160 0 1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1722_
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1723_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1724_
timestamp 1698431365
transform 1 0 12992 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1725_
timestamp 1698431365
transform -1 0 19152 0 1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1726_
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1727_
timestamp 1698431365
transform -1 0 41328 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1728_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41328 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1729_
timestamp 1698431365
transform 1 0 44464 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1730_
timestamp 1698431365
transform 1 0 39200 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1731_
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1732_
timestamp 1698431365
transform 1 0 33040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1733_
timestamp 1698431365
transform 1 0 30688 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1734_
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1735_
timestamp 1698431365
transform 1 0 27104 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1736_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1737_
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1738_
timestamp 1698431365
transform 1 0 29344 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1739_
timestamp 1698431365
transform 1 0 29568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform -1 0 32480 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1741_
timestamp 1698431365
transform -1 0 31920 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1742_
timestamp 1698431365
transform 1 0 19824 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1743_
timestamp 1698431365
transform 1 0 22512 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1744_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1745_
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1746_
timestamp 1698431365
transform -1 0 24192 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1747_
timestamp 1698431365
transform 1 0 22624 0 1 6272
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1748_
timestamp 1698431365
transform 1 0 30464 0 1 6272
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698431365
transform 1 0 40096 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1750_
timestamp 1698431365
transform 1 0 43792 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1751_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43568 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1752_
timestamp 1698431365
transform 1 0 45696 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1753_
timestamp 1698431365
transform -1 0 48944 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1754_
timestamp 1698431365
transform 1 0 46368 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1755_
timestamp 1698431365
transform 1 0 47040 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1756_
timestamp 1698431365
transform -1 0 48160 0 -1 4704
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1757_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1758_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1759_
timestamp 1698431365
transform -1 0 46480 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1760_
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1761_
timestamp 1698431365
transform -1 0 29792 0 -1 7840
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1762_
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1763_
timestamp 1698431365
transform 1 0 27440 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1764_
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1765_
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1766_
timestamp 1698431365
transform -1 0 24416 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1767_
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1768_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1769_
timestamp 1698431365
transform 1 0 27776 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1770_
timestamp 1698431365
transform 1 0 27216 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1771_
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1772_
timestamp 1698431365
transform 1 0 34944 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1773_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1774_
timestamp 1698431365
transform -1 0 29344 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1775_
timestamp 1698431365
transform -1 0 33040 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1776_
timestamp 1698431365
transform -1 0 31920 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1777_
timestamp 1698431365
transform 1 0 33936 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1778_
timestamp 1698431365
transform 1 0 33040 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1779_
timestamp 1698431365
transform 1 0 42448 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1780_
timestamp 1698431365
transform 1 0 42336 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1781_
timestamp 1698431365
transform -1 0 41552 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1782_
timestamp 1698431365
transform 1 0 43120 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1783_
timestamp 1698431365
transform 1 0 43008 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1784_
timestamp 1698431365
transform 1 0 44688 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1785_
timestamp 1698431365
transform -1 0 39312 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1786_
timestamp 1698431365
transform -1 0 37744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1787_
timestamp 1698431365
transform 1 0 21952 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1788_
timestamp 1698431365
transform 1 0 23744 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1789_
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1790_
timestamp 1698431365
transform 1 0 25984 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1791_
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1792_
timestamp 1698431365
transform 1 0 24976 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1793_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1794_
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1795_
timestamp 1698431365
transform 1 0 9632 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1796_
timestamp 1698431365
transform 1 0 25760 0 1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1797_
timestamp 1698431365
transform -1 0 29008 0 -1 12544
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1798_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1799_
timestamp 1698431365
transform -1 0 40432 0 -1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1800_
timestamp 1698431365
transform -1 0 22176 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1801_
timestamp 1698431365
transform -1 0 21952 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1698431365
transform -1 0 21728 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1803_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1804_
timestamp 1698431365
transform -1 0 23184 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1805_
timestamp 1698431365
transform -1 0 24752 0 -1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1806_
timestamp 1698431365
transform 1 0 19488 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1807_
timestamp 1698431365
transform 1 0 22848 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1808_
timestamp 1698431365
transform -1 0 25984 0 1 10976
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1809_
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1810_
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1811_
timestamp 1698431365
transform 1 0 42672 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1812_
timestamp 1698431365
transform 1 0 46144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1813_
timestamp 1698431365
transform 1 0 42000 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1814_
timestamp 1698431365
transform 1 0 46592 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1815_
timestamp 1698431365
transform -1 0 47824 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1816_
timestamp 1698431365
transform 1 0 44912 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1817_
timestamp 1698431365
transform 1 0 47040 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1818_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46480 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1819_
timestamp 1698431365
transform 1 0 46368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1820_
timestamp 1698431365
transform 1 0 46704 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1821_
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1822_
timestamp 1698431365
transform 1 0 47488 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1823_
timestamp 1698431365
transform 1 0 50176 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1824_
timestamp 1698431365
transform 1 0 51520 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1825_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43008 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1826_
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1827_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1828_
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1829_
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1830_
timestamp 1698431365
transform 1 0 12992 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1831_
timestamp 1698431365
transform 1 0 24192 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1832_
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1833_
timestamp 1698431365
transform -1 0 30800 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1834_
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1835_
timestamp 1698431365
transform -1 0 32704 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1836_
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1837_
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1838_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1839_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 17248
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1840_
timestamp 1698431365
transform 1 0 42672 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1841_
timestamp 1698431365
transform 1 0 45248 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1842_
timestamp 1698431365
transform 1 0 35056 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 38080 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1844_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1845_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28448 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1846_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26880 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1847_
timestamp 1698431365
transform 1 0 26992 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1848_
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1849_
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1850_
timestamp 1698431365
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1851_
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1852_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1853_
timestamp 1698431365
transform 1 0 33152 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1854_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1855_
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1856_
timestamp 1698431365
transform -1 0 37408 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform 1 0 39200 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1858_
timestamp 1698431365
transform -1 0 39424 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1859_
timestamp 1698431365
transform 1 0 22624 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1860_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29680 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1861_
timestamp 1698431365
transform 1 0 33040 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1862_
timestamp 1698431365
transform -1 0 34720 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1863_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1864_
timestamp 1698431365
transform -1 0 22624 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1866_
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1867_
timestamp 1698431365
transform 1 0 33488 0 -1 14112
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1868_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1869_
timestamp 1698431365
transform -1 0 26768 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _1870_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform -1 0 25760 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1872_
timestamp 1698431365
transform -1 0 22624 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1873_
timestamp 1698431365
transform 1 0 22400 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_4  _1874_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1875_
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1876_
timestamp 1698431365
transform -1 0 22624 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1877_
timestamp 1698431365
transform -1 0 26768 0 1 15680
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1878_
timestamp 1698431365
transform 1 0 37968 0 1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1879_
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1880_
timestamp 1698431365
transform 1 0 46592 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1881_
timestamp 1698431365
transform 1 0 46704 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1882_
timestamp 1698431365
transform 1 0 48944 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1698431365
transform 1 0 49280 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1884_
timestamp 1698431365
transform 1 0 50064 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1885_
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1886_
timestamp 1698431365
transform 1 0 47712 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1887_
timestamp 1698431365
transform 1 0 50400 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1888_
timestamp 1698431365
transform -1 0 50512 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1889_
timestamp 1698431365
transform 1 0 51520 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1890_
timestamp 1698431365
transform 1 0 47488 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1891_
timestamp 1698431365
transform 1 0 48608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1892_
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1893_
timestamp 1698431365
transform -1 0 51856 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1894_
timestamp 1698431365
transform 1 0 52192 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1895_
timestamp 1698431365
transform 1 0 53536 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1896_
timestamp 1698431365
transform -1 0 50064 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1897_
timestamp 1698431365
transform 1 0 50848 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1898_
timestamp 1698431365
transform 1 0 26544 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1899_
timestamp 1698431365
transform 1 0 25648 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1900_
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1901_
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1698431365
transform 1 0 31584 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1903_
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1904_
timestamp 1698431365
transform 1 0 32144 0 1 10976
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1906_
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1907_
timestamp 1698431365
transform 1 0 36064 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1908_
timestamp 1698431365
transform 1 0 39424 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1909_
timestamp 1698431365
transform -1 0 14000 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1910_
timestamp 1698431365
transform -1 0 24528 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1911_
timestamp 1698431365
transform -1 0 24752 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1912_
timestamp 1698431365
transform -1 0 19600 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1913_
timestamp 1698431365
transform 1 0 13104 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1914_
timestamp 1698431365
transform -1 0 18368 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1915_
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1916_
timestamp 1698431365
transform 1 0 19264 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1917_
timestamp 1698431365
transform -1 0 23632 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1918_
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1919_
timestamp 1698431365
transform -1 0 39200 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1920_
timestamp 1698431365
transform 1 0 46032 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1921_
timestamp 1698431365
transform -1 0 48384 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1922_
timestamp 1698431365
transform -1 0 42896 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1923_
timestamp 1698431365
transform -1 0 45248 0 -1 12544
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1924_
timestamp 1698431365
transform 1 0 40880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1925_
timestamp 1698431365
transform -1 0 26432 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform 1 0 27216 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1927_
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1928_
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1929_
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1930_
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1931_
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1932_
timestamp 1698431365
transform -1 0 24528 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1933_
timestamp 1698431365
transform -1 0 23520 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1934_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1935_
timestamp 1698431365
transform 1 0 33040 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1936_
timestamp 1698431365
transform -1 0 42336 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1937_
timestamp 1698431365
transform -1 0 42896 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1938_
timestamp 1698431365
transform 1 0 48384 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1939_
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1940_
timestamp 1698431365
transform -1 0 52080 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1941_
timestamp 1698431365
transform 1 0 52640 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1942_
timestamp 1698431365
transform 1 0 53424 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1943_
timestamp 1698431365
transform 1 0 54096 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1944_
timestamp 1698431365
transform 1 0 55440 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1945_
timestamp 1698431365
transform -1 0 39536 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1946_
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1947_
timestamp 1698431365
transform 1 0 28896 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1948_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1949_
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1950_
timestamp 1698431365
transform -1 0 18368 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1951_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1952_
timestamp 1698431365
transform -1 0 22064 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1953_
timestamp 1698431365
transform -1 0 31136 0 1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1954_
timestamp 1698431365
transform 1 0 43680 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1955_
timestamp 1698431365
transform 1 0 46928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1956_
timestamp 1698431365
transform 1 0 35504 0 -1 10976
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1957_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1698431365
transform -1 0 22512 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1959_
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1960_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1961_
timestamp 1698431365
transform 1 0 28224 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1962_
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1963_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1964_
timestamp 1698431365
transform -1 0 38752 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1965_
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1966_
timestamp 1698431365
transform -1 0 43232 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1967_
timestamp 1698431365
transform 1 0 42896 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1968_
timestamp 1698431365
transform -1 0 33600 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1969_
timestamp 1698431365
transform -1 0 32592 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1970_
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1971_
timestamp 1698431365
transform 1 0 27440 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1972_
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1973_
timestamp 1698431365
transform 1 0 25648 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1974_
timestamp 1698431365
transform 1 0 26320 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1975_
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1976_
timestamp 1698431365
transform -1 0 27104 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1977_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1978_
timestamp 1698431365
transform 1 0 29792 0 1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1979_
timestamp 1698431365
transform -1 0 44688 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1980_
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1981_
timestamp 1698431365
transform 1 0 49952 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1982_
timestamp 1698431365
transform 1 0 48720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1983_
timestamp 1698431365
transform 1 0 49392 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1984_
timestamp 1698431365
transform 1 0 49616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1985_
timestamp 1698431365
transform -1 0 51408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1986_
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1987_
timestamp 1698431365
transform -1 0 52304 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1988_
timestamp 1698431365
transform -1 0 52416 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1989_
timestamp 1698431365
transform 1 0 52528 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1990_
timestamp 1698431365
transform 1 0 53088 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1991_
timestamp 1698431365
transform 1 0 54096 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1992_
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1993_
timestamp 1698431365
transform -1 0 34496 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1994_
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1995_
timestamp 1698431365
transform -1 0 32032 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1996_
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1997_
timestamp 1698431365
transform 1 0 19712 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1998_
timestamp 1698431365
transform -1 0 34720 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1999_
timestamp 1698431365
transform 1 0 35728 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2000_
timestamp 1698431365
transform -1 0 43120 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform -1 0 35168 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2002_
timestamp 1698431365
transform -1 0 33264 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2003_
timestamp 1698431365
transform 1 0 33600 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2004_
timestamp 1698431365
transform 1 0 27888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2005_
timestamp 1698431365
transform 1 0 31024 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2006_
timestamp 1698431365
transform -1 0 34048 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2007_
timestamp 1698431365
transform 1 0 34160 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2008_
timestamp 1698431365
transform 1 0 33152 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2009_
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2010_
timestamp 1698431365
transform 1 0 34832 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2011_
timestamp 1698431365
transform -1 0 42336 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2012_
timestamp 1698431365
transform 1 0 42112 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2013_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2014_
timestamp 1698431365
transform 1 0 45920 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2015_
timestamp 1698431365
transform -1 0 47152 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2016_
timestamp 1698431365
transform 1 0 33152 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2017_
timestamp 1698431365
transform -1 0 30128 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2018_
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2019_
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2020_
timestamp 1698431365
transform 1 0 37632 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2021_
timestamp 1698431365
transform 1 0 43680 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2022_
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2023_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48944 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2024_
timestamp 1698431365
transform 1 0 48832 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2025_
timestamp 1698431365
transform -1 0 51184 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2026_
timestamp 1698431365
transform 1 0 50400 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2027_
timestamp 1698431365
transform 1 0 51408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2028_
timestamp 1698431365
transform -1 0 53088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2029_
timestamp 1698431365
transform 1 0 54096 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2030_
timestamp 1698431365
transform 1 0 53984 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2031_
timestamp 1698431365
transform 1 0 54768 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2032_
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2033_
timestamp 1698431365
transform 1 0 35168 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2034_
timestamp 1698431365
transform -1 0 37744 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2035_
timestamp 1698431365
transform -1 0 34048 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2036_
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2037_
timestamp 1698431365
transform 1 0 22176 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2038_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24752 0 -1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2039_
timestamp 1698431365
transform 1 0 22848 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2040_
timestamp 1698431365
transform 1 0 34608 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2041_
timestamp 1698431365
transform -1 0 42448 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2042_
timestamp 1698431365
transform 1 0 45920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2043_
timestamp 1698431365
transform 1 0 46144 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2044_
timestamp 1698431365
transform 1 0 34944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2045_
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2046_
timestamp 1698431365
transform 1 0 30240 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2047_
timestamp 1698431365
transform -1 0 31360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2048_
timestamp 1698431365
transform -1 0 40768 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2049_
timestamp 1698431365
transform -1 0 40208 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2050_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39088 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2051_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2052_
timestamp 1698431365
transform -1 0 42224 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2053_
timestamp 1698431365
transform 1 0 46816 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2054_
timestamp 1698431365
transform 1 0 50176 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2055_
timestamp 1698431365
transform 1 0 49280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2056_
timestamp 1698431365
transform 1 0 50064 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2057_
timestamp 1698431365
transform 1 0 50848 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2058_
timestamp 1698431365
transform 1 0 52752 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2059_
timestamp 1698431365
transform 1 0 51184 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2060_
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2061_
timestamp 1698431365
transform 1 0 52976 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2062_
timestamp 1698431365
transform -1 0 52528 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2063_
timestamp 1698431365
transform -1 0 54656 0 1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2064_
timestamp 1698431365
transform -1 0 53984 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2065_
timestamp 1698431365
transform -1 0 56224 0 -1 18816
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2066_
timestamp 1698431365
transform 1 0 53312 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2067_
timestamp 1698431365
transform 1 0 54656 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2068_
timestamp 1698431365
transform -1 0 47936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2069_
timestamp 1698431365
transform -1 0 47040 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2070_
timestamp 1698431365
transform -1 0 47936 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2071_
timestamp 1698431365
transform 1 0 34160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2072_
timestamp 1698431365
transform -1 0 35952 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2073_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2074_
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2075_
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2076_
timestamp 1698431365
transform 1 0 35056 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2077_
timestamp 1698431365
transform -1 0 38864 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2078_
timestamp 1698431365
transform -1 0 23296 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2079_
timestamp 1698431365
transform 1 0 25200 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2080_
timestamp 1698431365
transform 1 0 25984 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2081_
timestamp 1698431365
transform -1 0 35728 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2082_
timestamp 1698431365
transform 1 0 41440 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2083_
timestamp 1698431365
transform 1 0 41552 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698431365
transform 1 0 46816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2085_
timestamp 1698431365
transform 1 0 47600 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2086_
timestamp 1698431365
transform 1 0 49504 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2087_
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2088_
timestamp 1698431365
transform 1 0 31136 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2089_
timestamp 1698431365
transform 1 0 31360 0 1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2090_
timestamp 1698431365
transform 1 0 43008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2091_
timestamp 1698431365
transform 1 0 42784 0 -1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2092_
timestamp 1698431365
transform 1 0 49056 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2093_
timestamp 1698431365
transform 1 0 50960 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2094_
timestamp 1698431365
transform 1 0 51520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2095_
timestamp 1698431365
transform 1 0 52752 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2096_
timestamp 1698431365
transform 1 0 54096 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2097_
timestamp 1698431365
transform 1 0 54208 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2098_
timestamp 1698431365
transform 1 0 53424 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2099_
timestamp 1698431365
transform 1 0 53312 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2100_
timestamp 1698431365
transform -1 0 54992 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2101_
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2102_
timestamp 1698431365
transform -1 0 41328 0 1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2103_
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2104_
timestamp 1698431365
transform -1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2105_
timestamp 1698431365
transform 1 0 33936 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2106_
timestamp 1698431365
transform -1 0 45920 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2107_
timestamp 1698431365
transform -1 0 46144 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2108_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2109_
timestamp 1698431365
transform 1 0 46032 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2110_
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2111_
timestamp 1698431365
transform -1 0 34160 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2112_
timestamp 1698431365
transform 1 0 43232 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2113_
timestamp 1698431365
transform 1 0 42336 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2114_
timestamp 1698431365
transform 1 0 42896 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2115_
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2116_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2117_
timestamp 1698431365
transform 1 0 49056 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2118_
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2119_
timestamp 1698431365
transform 1 0 50400 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2120_
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2121_
timestamp 1698431365
transform -1 0 53312 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2122_
timestamp 1698431365
transform 1 0 52640 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2123_
timestamp 1698431365
transform 1 0 53200 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2124_
timestamp 1698431365
transform 1 0 54544 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2125_
timestamp 1698431365
transform 1 0 46816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2126_
timestamp 1698431365
transform 1 0 46928 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2127_
timestamp 1698431365
transform 1 0 48608 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2128_
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2129_
timestamp 1698431365
transform 1 0 34944 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2130_
timestamp 1698431365
transform 1 0 43120 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2131_
timestamp 1698431365
transform -1 0 43008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2132_
timestamp 1698431365
transform 1 0 45024 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2133_
timestamp 1698431365
transform -1 0 46928 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2134_
timestamp 1698431365
transform 1 0 45584 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2135_
timestamp 1698431365
transform -1 0 51296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2136_
timestamp 1698431365
transform 1 0 49280 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2137_
timestamp 1698431365
transform 1 0 51296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2138_
timestamp 1698431365
transform 1 0 50064 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2139_
timestamp 1698431365
transform -1 0 53424 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2140_
timestamp 1698431365
transform 1 0 52416 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2141_
timestamp 1698431365
transform 1 0 53760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2142_
timestamp 1698431365
transform -1 0 46816 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2143_
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2144_
timestamp 1698431365
transform 1 0 45696 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2145_
timestamp 1698431365
transform 1 0 49392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1698431365
transform -1 0 51968 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2147_
timestamp 1698431365
transform -1 0 53200 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2148_
timestamp 1698431365
transform -1 0 47376 0 1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2149_
timestamp 1698431365
transform 1 0 42336 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2150_
timestamp 1698431365
transform 1 0 43680 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2151_
timestamp 1698431365
transform -1 0 15008 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2152_
timestamp 1698431365
transform 1 0 14448 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2153_
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2154_
timestamp 1698431365
transform -1 0 19712 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2155_
timestamp 1698431365
transform 1 0 15008 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2156_
timestamp 1698431365
transform -1 0 19488 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2157_
timestamp 1698431365
transform 1 0 18032 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2158_
timestamp 1698431365
transform 1 0 22736 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2159_
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2160_
timestamp 1698431365
transform -1 0 22176 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2161_
timestamp 1698431365
transform -1 0 12768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2162_
timestamp 1698431365
transform 1 0 11536 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2163_
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2164_
timestamp 1698431365
transform -1 0 17024 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2165_
timestamp 1698431365
transform 1 0 18480 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2166_
timestamp 1698431365
transform 1 0 9968 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2167_
timestamp 1698431365
transform 1 0 9296 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2168_
timestamp 1698431365
transform -1 0 14224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2169_
timestamp 1698431365
transform 1 0 13552 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2170_
timestamp 1698431365
transform -1 0 27664 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2171_
timestamp 1698431365
transform -1 0 24864 0 -1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2172_
timestamp 1698431365
transform 1 0 29680 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2173_
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2174_
timestamp 1698431365
transform 1 0 9296 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2175_
timestamp 1698431365
transform 1 0 8624 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2176_
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2177_
timestamp 1698431365
transform -1 0 13104 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _2178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15904 0 1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2179_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2180_
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2181_
timestamp 1698431365
transform -1 0 13552 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2182_
timestamp 1698431365
transform 1 0 20832 0 -1 40768
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2183_
timestamp 1698431365
transform 1 0 26768 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2184_
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2185_
timestamp 1698431365
transform 1 0 29120 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2186_
timestamp 1698431365
transform -1 0 30016 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2187_
timestamp 1698431365
transform 1 0 27776 0 -1 40768
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2188_
timestamp 1698431365
transform -1 0 13776 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2189_
timestamp 1698431365
transform -1 0 16800 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2190_
timestamp 1698431365
transform 1 0 9856 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2191_
timestamp 1698431365
transform 1 0 11536 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2192_
timestamp 1698431365
transform 1 0 16352 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2193_
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2194_
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2195_
timestamp 1698431365
transform -1 0 18368 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2196_
timestamp 1698431365
transform -1 0 18368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2197_
timestamp 1698431365
transform -1 0 19712 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _2198_
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2199_
timestamp 1698431365
transform -1 0 27888 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2200_
timestamp 1698431365
transform -1 0 23520 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2201_
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2202_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2203_
timestamp 1698431365
transform 1 0 38640 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2204_
timestamp 1698431365
transform -1 0 44800 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2205_
timestamp 1698431365
transform 1 0 41440 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2206_
timestamp 1698431365
transform 1 0 42224 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2207_
timestamp 1698431365
transform -1 0 42448 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2208_
timestamp 1698431365
transform 1 0 30688 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2209_
timestamp 1698431365
transform 1 0 17808 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2210_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2211_
timestamp 1698431365
transform 1 0 14448 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2212_
timestamp 1698431365
transform 1 0 15456 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2213_
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2214_
timestamp 1698431365
transform 1 0 23856 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2215_
timestamp 1698431365
transform -1 0 27440 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2216_
timestamp 1698431365
transform 1 0 9856 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2217_
timestamp 1698431365
transform -1 0 20160 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2218_
timestamp 1698431365
transform -1 0 29904 0 -1 39200
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2219_
timestamp 1698431365
transform -1 0 14784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2220_
timestamp 1698431365
transform 1 0 11536 0 -1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2221_
timestamp 1698431365
transform 1 0 30912 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2222_
timestamp 1698431365
transform 1 0 29904 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2223_
timestamp 1698431365
transform 1 0 10640 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2224_
timestamp 1698431365
transform 1 0 14672 0 1 39200
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2225_
timestamp 1698431365
transform -1 0 15456 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2226_
timestamp 1698431365
transform -1 0 24416 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2227_
timestamp 1698431365
transform -1 0 24192 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2228_
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _2229_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31024 0 1 39200
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2230_
timestamp 1698431365
transform -1 0 40208 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2231_
timestamp 1698431365
transform 1 0 19376 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2232_
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2233_
timestamp 1698431365
transform 1 0 25648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2234_
timestamp 1698431365
transform -1 0 23632 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2235_
timestamp 1698431365
transform 1 0 9296 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2236_
timestamp 1698431365
transform 1 0 25760 0 -1 34496
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2237_
timestamp 1698431365
transform -1 0 14672 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2238_
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2239_
timestamp 1698431365
transform -1 0 30352 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2240_
timestamp 1698431365
transform 1 0 33488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2241_
timestamp 1698431365
transform 1 0 41776 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2242_
timestamp 1698431365
transform 1 0 42336 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2243_
timestamp 1698431365
transform 1 0 43344 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2244_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2245_
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2246_
timestamp 1698431365
transform -1 0 30800 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2247_
timestamp 1698431365
transform -1 0 23408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2248_
timestamp 1698431365
transform 1 0 17920 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2249_
timestamp 1698431365
transform -1 0 11200 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2250_
timestamp 1698431365
transform 1 0 10192 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2251_
timestamp 1698431365
transform 1 0 15344 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2252_
timestamp 1698431365
transform 1 0 18592 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2253_
timestamp 1698431365
transform 1 0 19152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2254_
timestamp 1698431365
transform -1 0 27216 0 -1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2255_
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2256_
timestamp 1698431365
transform 1 0 11312 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2257_
timestamp 1698431365
transform -1 0 19152 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2258_
timestamp 1698431365
transform -1 0 17920 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2259_
timestamp 1698431365
transform -1 0 10304 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2260_
timestamp 1698431365
transform 1 0 7168 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _2261_
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2262_
timestamp 1698431365
transform 1 0 24192 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2263_
timestamp 1698431365
transform -1 0 24528 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2264_
timestamp 1698431365
transform 1 0 25088 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2265_
timestamp 1698431365
transform -1 0 13104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2266_
timestamp 1698431365
transform -1 0 16016 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2267_
timestamp 1698431365
transform 1 0 27664 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2268_
timestamp 1698431365
transform -1 0 24752 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2269_
timestamp 1698431365
transform -1 0 23968 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2270_
timestamp 1698431365
transform -1 0 30464 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2271_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2272_
timestamp 1698431365
transform 1 0 38416 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2273_
timestamp 1698431365
transform 1 0 41328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2274_
timestamp 1698431365
transform -1 0 41328 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2275_
timestamp 1698431365
transform -1 0 22512 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2276_
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2277_
timestamp 1698431365
transform -1 0 24864 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2278_
timestamp 1698431365
transform 1 0 14672 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2279_
timestamp 1698431365
transform 1 0 12208 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2280_
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2281_
timestamp 1698431365
transform 1 0 23072 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2282_
timestamp 1698431365
transform 1 0 25088 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1698431365
transform 1 0 23520 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2284_
timestamp 1698431365
transform -1 0 26544 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2285_
timestamp 1698431365
transform 1 0 18592 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2286_
timestamp 1698431365
transform -1 0 15904 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2287_
timestamp 1698431365
transform 1 0 29120 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2288_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2289_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2290_
timestamp 1698431365
transform 1 0 33376 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2291_
timestamp 1698431365
transform -1 0 33712 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2292_
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2293_
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2294_
timestamp 1698431365
transform -1 0 35392 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2295_
timestamp 1698431365
transform 1 0 34384 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2296_
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2297_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2298_
timestamp 1698431365
transform 1 0 9520 0 -1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2299_
timestamp 1698431365
transform 1 0 13216 0 -1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _2300_
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2301_
timestamp 1698431365
transform 1 0 29120 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2302_
timestamp 1698431365
transform 1 0 30352 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2303_
timestamp 1698431365
transform 1 0 30912 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2304_
timestamp 1698431365
transform -1 0 35840 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2305_
timestamp 1698431365
transform 1 0 35840 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2306_
timestamp 1698431365
transform -1 0 39200 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2307_
timestamp 1698431365
transform 1 0 39200 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2308_
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2309_
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2310_
timestamp 1698431365
transform 1 0 43568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2311_
timestamp 1698431365
transform 1 0 46704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1698431365
transform 1 0 39088 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2313_
timestamp 1698431365
transform -1 0 40320 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2314_
timestamp 1698431365
transform -1 0 42224 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2315_
timestamp 1698431365
transform 1 0 38640 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2316_
timestamp 1698431365
transform 1 0 39872 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2317_
timestamp 1698431365
transform -1 0 22400 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2318_
timestamp 1698431365
transform -1 0 19040 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2319_
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2320_
timestamp 1698431365
transform 1 0 16128 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2321_
timestamp 1698431365
transform 1 0 12208 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2322_
timestamp 1698431365
transform 1 0 10416 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2323_
timestamp 1698431365
transform -1 0 27888 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2324_
timestamp 1698431365
transform -1 0 20832 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2325_
timestamp 1698431365
transform -1 0 19488 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2326_
timestamp 1698431365
transform 1 0 19488 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2327_
timestamp 1698431365
transform 1 0 31248 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2328_
timestamp 1698431365
transform 1 0 10864 0 -1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2329_
timestamp 1698431365
transform -1 0 19712 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2330_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2331_
timestamp 1698431365
transform -1 0 18368 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2332_
timestamp 1698431365
transform -1 0 27776 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2333_
timestamp 1698431365
transform -1 0 28224 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2334_
timestamp 1698431365
transform -1 0 32704 0 -1 42336
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2335_
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2336_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2337_
timestamp 1698431365
transform 1 0 33152 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2338_
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2339_
timestamp 1698431365
transform -1 0 26656 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2340_
timestamp 1698431365
transform -1 0 27216 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2341_
timestamp 1698431365
transform 1 0 18704 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2342_
timestamp 1698431365
transform 1 0 19488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2343_
timestamp 1698431365
transform 1 0 13440 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2344_
timestamp 1698431365
transform -1 0 9184 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2345_
timestamp 1698431365
transform -1 0 15456 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2346_
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2347_
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2348_
timestamp 1698431365
transform 1 0 25760 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2349_
timestamp 1698431365
transform 1 0 33600 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2350_
timestamp 1698431365
transform -1 0 36064 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2351_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2352_
timestamp 1698431365
transform 1 0 19152 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2353_
timestamp 1698431365
transform -1 0 17920 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2354_
timestamp 1698431365
transform 1 0 20832 0 -1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2355_
timestamp 1698431365
transform 1 0 17360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2356_
timestamp 1698431365
transform -1 0 15008 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2357_
timestamp 1698431365
transform 1 0 18256 0 -1 36064
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2358_
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2359_
timestamp 1698431365
transform 1 0 30912 0 1 36064
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2360_
timestamp 1698431365
transform 1 0 34608 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2361_
timestamp 1698431365
transform -1 0 34608 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2362_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2363_
timestamp 1698431365
transform 1 0 36064 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2364_
timestamp 1698431365
transform 1 0 43008 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2365_
timestamp 1698431365
transform 1 0 43344 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2366_
timestamp 1698431365
transform -1 0 43904 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2367_
timestamp 1698431365
transform 1 0 46592 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2368_
timestamp 1698431365
transform 1 0 46480 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2369_
timestamp 1698431365
transform 1 0 49056 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2370_
timestamp 1698431365
transform -1 0 46704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2371_
timestamp 1698431365
transform 1 0 46256 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2372_
timestamp 1698431365
transform 1 0 46704 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2373_
timestamp 1698431365
transform 1 0 35280 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2374_
timestamp 1698431365
transform -1 0 37744 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2375_
timestamp 1698431365
transform 1 0 45024 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2376_
timestamp 1698431365
transform -1 0 39760 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2377_
timestamp 1698431365
transform 1 0 39424 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2378_
timestamp 1698431365
transform -1 0 26208 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2379_
timestamp 1698431365
transform -1 0 23184 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2380_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2381_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2382_
timestamp 1698431365
transform -1 0 20944 0 1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2383_
timestamp 1698431365
transform -1 0 29344 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2384_
timestamp 1698431365
transform -1 0 17920 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2385_
timestamp 1698431365
transform -1 0 16800 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2386_
timestamp 1698431365
transform 1 0 19712 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2387_
timestamp 1698431365
transform -1 0 24864 0 -1 43904
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2388_
timestamp 1698431365
transform 1 0 41552 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2389_
timestamp 1698431365
transform 1 0 42896 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2390_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2391_
timestamp 1698431365
transform 1 0 41216 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2392_
timestamp 1698431365
transform 1 0 42672 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2393_
timestamp 1698431365
transform -1 0 45472 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2394_
timestamp 1698431365
transform 1 0 12544 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2395_
timestamp 1698431365
transform 1 0 16464 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2396_
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2397_
timestamp 1698431365
transform -1 0 16352 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2398_
timestamp 1698431365
transform 1 0 25200 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2399_
timestamp 1698431365
transform -1 0 16352 0 1 42336
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2400_
timestamp 1698431365
transform 1 0 14560 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2401_
timestamp 1698431365
transform 1 0 21168 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2402_
timestamp 1698431365
transform 1 0 21728 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2403_
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2404_
timestamp 1698431365
transform 1 0 11648 0 -1 45472
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2405_
timestamp 1698431365
transform 1 0 21616 0 1 45472
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2406_
timestamp 1698431365
transform 1 0 34832 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2407_
timestamp 1698431365
transform 1 0 34496 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2408_
timestamp 1698431365
transform -1 0 21840 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2409_
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2410_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2411_
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2412_
timestamp 1698431365
transform -1 0 20720 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2413_
timestamp 1698431365
transform 1 0 19712 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2414_
timestamp 1698431365
transform 1 0 20160 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2415_
timestamp 1698431365
transform 1 0 10640 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2416_
timestamp 1698431365
transform -1 0 24864 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2417_
timestamp 1698431365
transform -1 0 14784 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2418_
timestamp 1698431365
transform 1 0 22960 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2419_
timestamp 1698431365
transform 1 0 25760 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2420_
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2421_
timestamp 1698431365
transform 1 0 24752 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2422_
timestamp 1698431365
transform -1 0 25760 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2423_
timestamp 1698431365
transform 1 0 31472 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2424_
timestamp 1698431365
transform 1 0 34832 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2425_
timestamp 1698431365
transform 1 0 33488 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2426_
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2427_
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2428_
timestamp 1698431365
transform 1 0 45696 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2429_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2430_
timestamp 1698431365
transform 1 0 49952 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2431_
timestamp 1698431365
transform -1 0 27664 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2432_
timestamp 1698431365
transform -1 0 27776 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2433_
timestamp 1698431365
transform 1 0 13552 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2434_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26880 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2435_
timestamp 1698431365
transform 1 0 27888 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2436_
timestamp 1698431365
transform 1 0 27888 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2437_
timestamp 1698431365
transform 1 0 13104 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2438_
timestamp 1698431365
transform 1 0 23744 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2439_
timestamp 1698431365
transform 1 0 26544 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2440_
timestamp 1698431365
transform 1 0 17696 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2441_
timestamp 1698431365
transform 1 0 27104 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2442_
timestamp 1698431365
transform 1 0 14448 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2443_
timestamp 1698431365
transform 1 0 15120 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2444_
timestamp 1698431365
transform -1 0 30240 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2445_
timestamp 1698431365
transform -1 0 39424 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2446_
timestamp 1698431365
transform 1 0 37744 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2447_
timestamp 1698431365
transform 1 0 38304 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2448_
timestamp 1698431365
transform -1 0 43680 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2449_
timestamp 1698431365
transform 1 0 42112 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2450_
timestamp 1698431365
transform 1 0 34048 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1698431365
transform 1 0 35840 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2452_
timestamp 1698431365
transform -1 0 14224 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2453_
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2454_
timestamp 1698431365
transform 1 0 14784 0 1 48608
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2455_
timestamp 1698431365
transform 1 0 18144 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2456_
timestamp 1698431365
transform 1 0 19264 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1698431365
transform -1 0 23408 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2458_
timestamp 1698431365
transform 1 0 16464 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2459_
timestamp 1698431365
transform 1 0 17584 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform -1 0 20944 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2461_
timestamp 1698431365
transform -1 0 19040 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2462_
timestamp 1698431365
transform -1 0 19488 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1698431365
transform 1 0 18704 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2464_
timestamp 1698431365
transform -1 0 22960 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2465_
timestamp 1698431365
transform 1 0 37632 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2466_
timestamp 1698431365
transform -1 0 38080 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _2467_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33488 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2468_
timestamp 1698431365
transform 1 0 34160 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2469_
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2470_
timestamp 1698431365
transform 1 0 17136 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2471_
timestamp 1698431365
transform -1 0 27104 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2472_
timestamp 1698431365
transform 1 0 27440 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2473_
timestamp 1698431365
transform -1 0 32032 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2474_
timestamp 1698431365
transform 1 0 34160 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2475_
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2476_
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2477_
timestamp 1698431365
transform 1 0 47040 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2478_
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2479_
timestamp 1698431365
transform 1 0 44352 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2480_
timestamp 1698431365
transform 1 0 45248 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2481_
timestamp 1698431365
transform 1 0 46480 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2482_
timestamp 1698431365
transform 1 0 48944 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2483_
timestamp 1698431365
transform 1 0 45248 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2484_
timestamp 1698431365
transform 1 0 46144 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2485_
timestamp 1698431365
transform 1 0 48384 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2486_
timestamp 1698431365
transform 1 0 49952 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2487_
timestamp 1698431365
transform 1 0 51296 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2488_
timestamp 1698431365
transform 1 0 46144 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2489_
timestamp 1698431365
transform -1 0 47824 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2490_
timestamp 1698431365
transform 1 0 44016 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2491_
timestamp 1698431365
transform -1 0 11984 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2492_
timestamp 1698431365
transform -1 0 31024 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2493_
timestamp 1698431365
transform -1 0 26544 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2494_
timestamp 1698431365
transform -1 0 17472 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2495_
timestamp 1698431365
transform -1 0 22064 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2496_
timestamp 1698431365
transform 1 0 18368 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2497_
timestamp 1698431365
transform 1 0 11760 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2498_
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2499_
timestamp 1698431365
transform -1 0 14336 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform 1 0 20384 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2501_
timestamp 1698431365
transform 1 0 22848 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2502_
timestamp 1698431365
transform -1 0 23296 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2503_
timestamp 1698431365
transform 1 0 23408 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2504_
timestamp 1698431365
transform -1 0 39760 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2505_
timestamp 1698431365
transform 1 0 43568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2506_
timestamp 1698431365
transform 1 0 34048 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2507_
timestamp 1698431365
transform 1 0 36064 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2508_
timestamp 1698431365
transform -1 0 31472 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2509_
timestamp 1698431365
transform -1 0 27888 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2510_
timestamp 1698431365
transform -1 0 23744 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2511_
timestamp 1698431365
transform 1 0 23520 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2513_
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2514_
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1698431365
transform 1 0 45360 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2516_
timestamp 1698431365
transform 1 0 11312 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2517_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2518_
timestamp 1698431365
transform 1 0 22176 0 1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2519_
timestamp 1698431365
transform -1 0 31584 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2520_
timestamp 1698431365
transform 1 0 30464 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2521_
timestamp 1698431365
transform -1 0 30352 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2522_
timestamp 1698431365
transform 1 0 29568 0 1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2523_
timestamp 1698431365
transform -1 0 34944 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2524_
timestamp 1698431365
transform 1 0 34720 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2525_
timestamp 1698431365
transform 1 0 44912 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2526_
timestamp 1698431365
transform 1 0 45808 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2527_
timestamp 1698431365
transform 1 0 49392 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2528_
timestamp 1698431365
transform 1 0 49392 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2529_
timestamp 1698431365
transform 1 0 50736 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2530_
timestamp 1698431365
transform 1 0 49392 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2531_
timestamp 1698431365
transform 1 0 50288 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2532_
timestamp 1698431365
transform 1 0 51968 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2533_
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2534_
timestamp 1698431365
transform -1 0 40320 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2535_
timestamp 1698431365
transform -1 0 38752 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2536_
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2537_
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2538_
timestamp 1698431365
transform 1 0 23632 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2539_
timestamp 1698431365
transform 1 0 14672 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2540_
timestamp 1698431365
transform -1 0 17024 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2541_
timestamp 1698431365
transform -1 0 16912 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2542_
timestamp 1698431365
transform 1 0 14448 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2543_
timestamp 1698431365
transform -1 0 22848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2544_
timestamp 1698431365
transform -1 0 23184 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2545_
timestamp 1698431365
transform 1 0 24080 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2546_
timestamp 1698431365
transform 1 0 23184 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2547_
timestamp 1698431365
transform -1 0 24304 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2548_
timestamp 1698431365
transform 1 0 39088 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2549_
timestamp 1698431365
transform -1 0 45248 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2550_
timestamp 1698431365
transform -1 0 33936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2551_
timestamp 1698431365
transform -1 0 34720 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2552_
timestamp 1698431365
transform -1 0 33600 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2553_
timestamp 1698431365
transform 1 0 17360 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2554_
timestamp 1698431365
transform 1 0 16576 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2555_
timestamp 1698431365
transform 1 0 15568 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2556_
timestamp 1698431365
transform -1 0 20048 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2557_
timestamp 1698431365
transform -1 0 17808 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2558_
timestamp 1698431365
transform 1 0 15344 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2559_
timestamp 1698431365
transform 1 0 30464 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2560_
timestamp 1698431365
transform 1 0 33600 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2561_
timestamp 1698431365
transform 1 0 42896 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2562_
timestamp 1698431365
transform -1 0 19936 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2563_
timestamp 1698431365
transform -1 0 30688 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2564_
timestamp 1698431365
transform -1 0 22064 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2565_
timestamp 1698431365
transform 1 0 19264 0 -1 54880
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2566_
timestamp 1698431365
transform 1 0 25424 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2567_
timestamp 1698431365
transform -1 0 21616 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2568_
timestamp 1698431365
transform -1 0 37744 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2569_
timestamp 1698431365
transform -1 0 35728 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2570_
timestamp 1698431365
transform -1 0 38304 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2571_
timestamp 1698431365
transform -1 0 50736 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2572_
timestamp 1698431365
transform 1 0 49504 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2573_
timestamp 1698431365
transform 1 0 45248 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2574_
timestamp 1698431365
transform -1 0 47152 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2575_
timestamp 1698431365
transform 1 0 46480 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2576_
timestamp 1698431365
transform 1 0 50064 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2577_
timestamp 1698431365
transform 1 0 50064 0 -1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2578_
timestamp 1698431365
transform 1 0 51184 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2579_
timestamp 1698431365
transform -1 0 54208 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2580_
timestamp 1698431365
transform 1 0 52640 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2581_
timestamp 1698431365
transform 1 0 49728 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2582_
timestamp 1698431365
transform 1 0 48832 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2583_
timestamp 1698431365
transform 1 0 50736 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2584_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2585_
timestamp 1698431365
transform -1 0 44016 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2586_
timestamp 1698431365
transform -1 0 41552 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2587_
timestamp 1698431365
transform 1 0 22288 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2588_
timestamp 1698431365
transform 1 0 27664 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2589_
timestamp 1698431365
transform 1 0 23296 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2590_
timestamp 1698431365
transform 1 0 23632 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2591_
timestamp 1698431365
transform 1 0 26656 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2592_
timestamp 1698431365
transform -1 0 30016 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2593_
timestamp 1698431365
transform 1 0 28000 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2594_
timestamp 1698431365
transform 1 0 27440 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2595_
timestamp 1698431365
transform -1 0 23632 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2596_
timestamp 1698431365
transform 1 0 24416 0 1 51744
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2597_
timestamp 1698431365
transform 1 0 26544 0 1 51744
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2598_
timestamp 1698431365
transform 1 0 39424 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2599_
timestamp 1698431365
transform 1 0 37408 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2600_
timestamp 1698431365
transform -1 0 39536 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2601_
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2602_
timestamp 1698431365
transform 1 0 42000 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2603_
timestamp 1698431365
transform 1 0 23632 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2604_
timestamp 1698431365
transform -1 0 25648 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2605_
timestamp 1698431365
transform 1 0 19712 0 1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2606_
timestamp 1698431365
transform -1 0 25984 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2607_
timestamp 1698431365
transform 1 0 35840 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2608_
timestamp 1698431365
transform 1 0 30688 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2609_
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2610_
timestamp 1698431365
transform -1 0 20384 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2611_
timestamp 1698431365
transform 1 0 19040 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2612_
timestamp 1698431365
transform 1 0 31584 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2613_
timestamp 1698431365
transform -1 0 36960 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2614_
timestamp 1698431365
transform 1 0 33936 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2615_
timestamp 1698431365
transform 1 0 33936 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2616_
timestamp 1698431365
transform 1 0 41440 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2617_
timestamp 1698431365
transform 1 0 42896 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2618_
timestamp 1698431365
transform -1 0 51968 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2619_
timestamp 1698431365
transform 1 0 51632 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2620_
timestamp 1698431365
transform -1 0 51744 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2621_
timestamp 1698431365
transform -1 0 53088 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2622_
timestamp 1698431365
transform 1 0 49168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2623_
timestamp 1698431365
transform 1 0 50624 0 -1 47040
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2624_
timestamp 1698431365
transform 1 0 51968 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2625_
timestamp 1698431365
transform 1 0 53424 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2626_
timestamp 1698431365
transform -1 0 40544 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2627_
timestamp 1698431365
transform 1 0 20384 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2628_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23072 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2629_
timestamp 1698431365
transform 1 0 15904 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2630_
timestamp 1698431365
transform 1 0 18928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2631_
timestamp 1698431365
transform 1 0 21728 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2632_
timestamp 1698431365
transform -1 0 23296 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2633_
timestamp 1698431365
transform -1 0 39760 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2634_
timestamp 1698431365
transform 1 0 40656 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2635_
timestamp 1698431365
transform 1 0 18928 0 -1 51744
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2636_
timestamp 1698431365
transform 1 0 33040 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2637_
timestamp 1698431365
transform 1 0 31696 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2638_
timestamp 1698431365
transform 1 0 35392 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2639_
timestamp 1698431365
transform 1 0 33936 0 1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2640_
timestamp 1698431365
transform 1 0 34160 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2641_
timestamp 1698431365
transform 1 0 25536 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2642_
timestamp 1698431365
transform 1 0 25536 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2643_
timestamp 1698431365
transform -1 0 27216 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2644_
timestamp 1698431365
transform 1 0 19488 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2645_
timestamp 1698431365
transform 1 0 24976 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2646_
timestamp 1698431365
transform 1 0 25648 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2647_
timestamp 1698431365
transform 1 0 26320 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2648_
timestamp 1698431365
transform -1 0 27552 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2649_
timestamp 1698431365
transform 1 0 31472 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2650_
timestamp 1698431365
transform 1 0 33264 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2651_
timestamp 1698431365
transform 1 0 33600 0 1 53312
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2652_
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2653_
timestamp 1698431365
transform 1 0 41104 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2654_
timestamp 1698431365
transform -1 0 44352 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2655_
timestamp 1698431365
transform 1 0 43120 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2656_
timestamp 1698431365
transform -1 0 51632 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2657_
timestamp 1698431365
transform 1 0 50512 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2658_
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2659_
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2660_
timestamp 1698431365
transform 1 0 41216 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2661_
timestamp 1698431365
transform 1 0 23072 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2662_
timestamp 1698431365
transform 1 0 24752 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2663_
timestamp 1698431365
transform 1 0 31024 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2664_
timestamp 1698431365
transform 1 0 30688 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2665_
timestamp 1698431365
transform -1 0 39760 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2666_
timestamp 1698431365
transform 1 0 39760 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2667_
timestamp 1698431365
transform -1 0 34496 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2668_
timestamp 1698431365
transform 1 0 33936 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2669_
timestamp 1698431365
transform 1 0 31136 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2670_
timestamp 1698431365
transform 1 0 32816 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2671_
timestamp 1698431365
transform -1 0 35168 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2672_
timestamp 1698431365
transform 1 0 27776 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2673_
timestamp 1698431365
transform 1 0 27776 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2674_
timestamp 1698431365
transform -1 0 31584 0 1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2675_
timestamp 1698431365
transform -1 0 34384 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2676_
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2677_
timestamp 1698431365
transform 1 0 38528 0 1 54880
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2678_
timestamp 1698431365
transform 1 0 41888 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2679_
timestamp 1698431365
transform 1 0 41888 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2680_
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2681_
timestamp 1698431365
transform 1 0 43456 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2682_
timestamp 1698431365
transform -1 0 50512 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2683_
timestamp 1698431365
transform 1 0 49616 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2684_
timestamp 1698431365
transform -1 0 52080 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2685_
timestamp 1698431365
transform 1 0 48944 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2686_
timestamp 1698431365
transform -1 0 52528 0 -1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2687_
timestamp 1698431365
transform 1 0 44576 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2688_
timestamp 1698431365
transform 1 0 45248 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2689_
timestamp 1698431365
transform 1 0 35728 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2690_
timestamp 1698431365
transform 1 0 27664 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2691_
timestamp 1698431365
transform 1 0 28672 0 -1 54880
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2692_
timestamp 1698431365
transform -1 0 35840 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2693_
timestamp 1698431365
transform 1 0 33712 0 -1 54880
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2694_
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2695_
timestamp 1698431365
transform -1 0 29904 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2696_
timestamp 1698431365
transform 1 0 29456 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2697_
timestamp 1698431365
transform 1 0 41664 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2698_
timestamp 1698431365
transform 1 0 42000 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2699_
timestamp 1698431365
transform 1 0 41776 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2700_
timestamp 1698431365
transform 1 0 43792 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2701_
timestamp 1698431365
transform 1 0 44912 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2702_
timestamp 1698431365
transform 1 0 37744 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2703_
timestamp 1698431365
transform 1 0 38640 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2704_
timestamp 1698431365
transform 1 0 38640 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2705_
timestamp 1698431365
transform 1 0 45584 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2706_
timestamp 1698431365
transform 1 0 47040 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2707_
timestamp 1698431365
transform 1 0 46592 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2708_
timestamp 1698431365
transform 1 0 47712 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2709_
timestamp 1698431365
transform 1 0 43904 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2710_
timestamp 1698431365
transform 1 0 45584 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2711_
timestamp 1698431365
transform 1 0 29120 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2712_
timestamp 1698431365
transform -1 0 31584 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2713_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38752 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2714_
timestamp 1698431365
transform 1 0 39200 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2715_
timestamp 1698431365
transform 1 0 45248 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2716_
timestamp 1698431365
transform 1 0 45584 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2717_
timestamp 1698431365
transform -1 0 47600 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2718_
timestamp 1698431365
transform 1 0 46480 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2719_
timestamp 1698431365
transform 1 0 47488 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2720_
timestamp 1698431365
transform 1 0 46032 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2721_
timestamp 1698431365
transform -1 0 47488 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2722_
timestamp 1698431365
transform 1 0 47488 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2723_
timestamp 1698431365
transform 1 0 48944 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2724_
timestamp 1698431365
transform 1 0 47040 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2725_
timestamp 1698431365
transform 1 0 43120 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2726_
timestamp 1698431365
transform 1 0 44912 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2727_
timestamp 1698431365
transform 1 0 45808 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2728_
timestamp 1698431365
transform 1 0 47152 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2729_
timestamp 1698431365
transform 1 0 47376 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2730_
timestamp 1698431365
transform -1 0 49056 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2731_
timestamp 1698431365
transform 1 0 45360 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2732_
timestamp 1698431365
transform 1 0 46256 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2733_
timestamp 1698431365
transform -1 0 43680 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2734_
timestamp 1698431365
transform -1 0 43120 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2735_
timestamp 1698431365
transform -1 0 26320 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2736_
timestamp 1698431365
transform 1 0 23072 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2737_
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2738_
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2739_
timestamp 1698431365
transform -1 0 23408 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2740_
timestamp 1698431365
transform -1 0 18480 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2741_
timestamp 1698431365
transform 1 0 18480 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2742_
timestamp 1698431365
transform 1 0 17584 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2743_
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2744_
timestamp 1698431365
transform 1 0 17920 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2745_
timestamp 1698431365
transform 1 0 23632 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2746_
timestamp 1698431365
transform -1 0 24192 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2747_
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2748_
timestamp 1698431365
transform 1 0 24192 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2749_
timestamp 1698431365
transform 1 0 24080 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2750_
timestamp 1698431365
transform 1 0 24192 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2751_
timestamp 1698431365
transform -1 0 24080 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2752_
timestamp 1698431365
transform 1 0 25312 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2753_
timestamp 1698431365
transform -1 0 25536 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2754_
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2755_
timestamp 1698431365
transform 1 0 26320 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2756_
timestamp 1698431365
transform -1 0 19040 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2757_
timestamp 1698431365
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2758_
timestamp 1698431365
transform 1 0 18256 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2759_
timestamp 1698431365
transform 1 0 18480 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2760_
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2761_
timestamp 1698431365
transform -1 0 20832 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2762_
timestamp 1698431365
transform -1 0 6720 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2763_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2764_
timestamp 1698431365
transform -1 0 22400 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2765_
timestamp 1698431365
transform -1 0 10192 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2766_
timestamp 1698431365
transform -1 0 25424 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2767_
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2768_
timestamp 1698431365
transform 1 0 22960 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2769_
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2770_
timestamp 1698431365
transform -1 0 23296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2771_
timestamp 1698431365
transform -1 0 12656 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2772_
timestamp 1698431365
transform -1 0 23744 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2773_
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2774_
timestamp 1698431365
transform -1 0 43680 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2775_
timestamp 1698431365
transform -1 0 43232 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2776_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41552 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2777_
timestamp 1698431365
transform 1 0 41328 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2778_
timestamp 1698431365
transform 1 0 29792 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2779_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2780_
timestamp 1698431365
transform 1 0 29568 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2781_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2782_
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2783_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2784_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2785_
timestamp 1698431365
transform -1 0 12880 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2786_
timestamp 1698431365
transform 1 0 5376 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2787_
timestamp 1698431365
transform -1 0 22848 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _2788_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2789_
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2790_
timestamp 1698431365
transform 1 0 34384 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2791_
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2792_
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_2  _2793_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4816 0 -1 25088
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2794_
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2795_
timestamp 1698431365
transform 1 0 5264 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_2  _2796_
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_2  _2797_
timestamp 1698431365
transform 1 0 11088 0 -1 26656
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2798_
timestamp 1698431365
transform -1 0 19040 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2799_
timestamp 1698431365
transform 1 0 34944 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2800_
timestamp 1698431365
transform 1 0 41552 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2801_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__I
timestamp 1698431365
transform -1 0 11424 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__I
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1393__I
timestamp 1698431365
transform 1 0 29344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__A1
timestamp 1698431365
transform 1 0 31136 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__I
timestamp 1698431365
transform 1 0 28672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A1
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform -1 0 32032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__B1
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__A2
timestamp 1698431365
transform 1 0 28560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__A4
timestamp 1698431365
transform 1 0 29232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__A1
timestamp 1698431365
transform 1 0 8400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1436__A1
timestamp 1698431365
transform 1 0 10416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__B
timestamp 1698431365
transform -1 0 12768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A1
timestamp 1698431365
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1698431365
transform 1 0 13216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__A2
timestamp 1698431365
transform -1 0 14000 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__A2
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A1
timestamp 1698431365
transform 1 0 35952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A2
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__I
timestamp 1698431365
transform 1 0 31696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__I
timestamp 1698431365
transform -1 0 34608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__I
timestamp 1698431365
transform 1 0 38080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__A1
timestamp 1698431365
transform -1 0 38864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A1
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1698431365
transform 1 0 36848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__A1
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A1
timestamp 1698431365
transform -1 0 26768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A2
timestamp 1698431365
transform -1 0 26992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__A2
timestamp 1698431365
transform 1 0 30800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__I
timestamp 1698431365
transform -1 0 10528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__I
timestamp 1698431365
transform 1 0 26096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__I
timestamp 1698431365
transform -1 0 23296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A2
timestamp 1698431365
transform -1 0 28448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__B
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__I
timestamp 1698431365
transform -1 0 6944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__B2
timestamp 1698431365
transform -1 0 27888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__C
timestamp 1698431365
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A1
timestamp 1698431365
transform -1 0 19040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A3
timestamp 1698431365
transform -1 0 16128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__I
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A1
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A2
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A1
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__I
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A1
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A1
timestamp 1698431365
transform -1 0 42896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A2
timestamp 1698431365
transform 1 0 11984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A2
timestamp 1698431365
transform -1 0 10752 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__I
timestamp 1698431365
transform -1 0 7840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A1
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A1
timestamp 1698431365
transform -1 0 9744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1698431365
transform -1 0 7392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A1
timestamp 1698431365
transform 1 0 6496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__I
timestamp 1698431365
transform -1 0 7616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A2
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A3
timestamp 1698431365
transform 1 0 8960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__B
timestamp 1698431365
transform -1 0 9632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A3
timestamp 1698431365
transform -1 0 6272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__A2
timestamp 1698431365
transform -1 0 5712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__A1
timestamp 1698431365
transform -1 0 10864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform -1 0 39200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1698431365
transform -1 0 6272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__A2
timestamp 1698431365
transform 1 0 10304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A2
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__I
timestamp 1698431365
transform 1 0 10528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A2
timestamp 1698431365
transform -1 0 8512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A1
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A2
timestamp 1698431365
transform -1 0 11200 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__B1
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__C
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I0
timestamp 1698431365
transform -1 0 8736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I1
timestamp 1698431365
transform 1 0 10640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__A1
timestamp 1698431365
transform -1 0 19600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__A2
timestamp 1698431365
transform -1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1698431365
transform 1 0 18480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A2
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__I
timestamp 1698431365
transform -1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__I
timestamp 1698431365
transform -1 0 10976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A1
timestamp 1698431365
transform -1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A1
timestamp 1698431365
transform -1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__I
timestamp 1698431365
transform 1 0 9856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A2
timestamp 1698431365
transform -1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A2
timestamp 1698431365
transform 1 0 11648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A1
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__I
timestamp 1698431365
transform 1 0 9744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A2
timestamp 1698431365
transform -1 0 12320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__B2
timestamp 1698431365
transform -1 0 13888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1698431365
transform -1 0 36624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A1
timestamp 1698431365
transform 1 0 37296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A1
timestamp 1698431365
transform -1 0 9408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A2
timestamp 1698431365
transform -1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A1
timestamp 1698431365
transform -1 0 15232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1698431365
transform -1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A1
timestamp 1698431365
transform -1 0 10192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__B
timestamp 1698431365
transform -1 0 16128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A1
timestamp 1698431365
transform 1 0 10080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__I0
timestamp 1698431365
transform -1 0 6720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A2
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A1
timestamp 1698431365
transform 1 0 9632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A2
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1698431365
transform 1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__B
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__A1
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A2
timestamp 1698431365
transform -1 0 17696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1698431365
transform 1 0 7168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__B
timestamp 1698431365
transform -1 0 6944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A1
timestamp 1698431365
transform -1 0 10752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1698431365
transform 1 0 6944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A2
timestamp 1698431365
transform -1 0 8512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__B
timestamp 1698431365
transform -1 0 8064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A2
timestamp 1698431365
transform -1 0 7840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__B
timestamp 1698431365
transform -1 0 8288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1698431365
transform -1 0 6496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__B
timestamp 1698431365
transform -1 0 6048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__B
timestamp 1698431365
transform -1 0 7392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A2
timestamp 1698431365
transform -1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A3
timestamp 1698431365
transform 1 0 39312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform 1 0 33152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A3
timestamp 1698431365
transform -1 0 30912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__B1
timestamp 1698431365
transform 1 0 33264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__B2
timestamp 1698431365
transform -1 0 29568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A3
timestamp 1698431365
transform -1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__I
timestamp 1698431365
transform 1 0 35728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__B
timestamp 1698431365
transform -1 0 31472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__I
timestamp 1698431365
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__I
timestamp 1698431365
transform 1 0 35056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1698431365
transform 1 0 34944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1698431365
transform 1 0 43456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1698431365
transform -1 0 43568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A2
timestamp 1698431365
transform -1 0 11312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__B
timestamp 1698431365
transform -1 0 11760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1698431365
transform 1 0 8736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__B
timestamp 1698431365
transform -1 0 11424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A1
timestamp 1698431365
transform -1 0 9296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A2
timestamp 1698431365
transform 1 0 9744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__B
timestamp 1698431365
transform -1 0 10416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A1
timestamp 1698431365
transform -1 0 11872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__B
timestamp 1698431365
transform -1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A2
timestamp 1698431365
transform 1 0 35952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__A1
timestamp 1698431365
transform 1 0 38416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A1
timestamp 1698431365
transform 1 0 36848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__B
timestamp 1698431365
transform -1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A1
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__B
timestamp 1698431365
transform -1 0 8960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1698431365
transform -1 0 6160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__B2
timestamp 1698431365
transform -1 0 9968 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A1
timestamp 1698431365
transform -1 0 8064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__B
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A1
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A1
timestamp 1698431365
transform 1 0 42336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A2
timestamp 1698431365
transform 1 0 40208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__A2
timestamp 1698431365
transform -1 0 41328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__B
timestamp 1698431365
transform -1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A2
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__I
timestamp 1698431365
transform 1 0 35168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A2
timestamp 1698431365
transform -1 0 30016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__B
timestamp 1698431365
transform -1 0 30464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__I
timestamp 1698431365
transform 1 0 34496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A1
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A2
timestamp 1698431365
transform -1 0 20384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__I
timestamp 1698431365
transform 1 0 33600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1698431365
transform 1 0 32144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1698431365
transform 1 0 33712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A1
timestamp 1698431365
transform -1 0 29120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__B
timestamp 1698431365
transform -1 0 31360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A2
timestamp 1698431365
transform -1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A2
timestamp 1698431365
transform -1 0 34272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__B1
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__C
timestamp 1698431365
transform -1 0 14896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1698431365
transform -1 0 35168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1698431365
transform 1 0 45584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__B
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A1
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__I
timestamp 1698431365
transform -1 0 27440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__A2
timestamp 1698431365
transform -1 0 17808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A2
timestamp 1698431365
transform 1 0 15232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698431365
transform -1 0 20608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1698431365
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A1
timestamp 1698431365
transform -1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__I
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1698431365
transform -1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A1
timestamp 1698431365
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__B
timestamp 1698431365
transform -1 0 34384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__A1
timestamp 1698431365
transform 1 0 45808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__I
timestamp 1698431365
transform 1 0 39536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__A1
timestamp 1698431365
transform 1 0 38416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1698431365
transform -1 0 19936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1698431365
transform -1 0 21392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__B
timestamp 1698431365
transform -1 0 21840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__I
timestamp 1698431365
transform -1 0 18928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__B
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A2
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__B
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A1
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A2
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A3
timestamp 1698431365
transform -1 0 38528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__B
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A1
timestamp 1698431365
transform 1 0 14112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A1
timestamp 1698431365
transform 1 0 21728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__B
timestamp 1698431365
transform 1 0 21280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__B
timestamp 1698431365
transform 1 0 19712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__I
timestamp 1698431365
transform -1 0 19488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__B
timestamp 1698431365
transform 1 0 45920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A2
timestamp 1698431365
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A1
timestamp 1698431365
transform 1 0 27104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A2
timestamp 1698431365
transform 1 0 31024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A2
timestamp 1698431365
transform -1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1698431365
transform 1 0 28112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A3
timestamp 1698431365
transform -1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A2
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 46368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A1
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A2
timestamp 1698431365
transform 1 0 35616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A3
timestamp 1698431365
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A2
timestamp 1698431365
transform -1 0 19488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__B2
timestamp 1698431365
transform 1 0 35392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__B
timestamp 1698431365
transform 1 0 34048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1698431365
transform -1 0 27664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__I
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A3
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__C
timestamp 1698431365
transform 1 0 35280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A1
timestamp 1698431365
transform -1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A2
timestamp 1698431365
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__B
timestamp 1698431365
transform -1 0 35952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__B2
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A1
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A2
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__B
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A3
timestamp 1698431365
transform -1 0 15680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__A1
timestamp 1698431365
transform -1 0 35168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__B2
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A2
timestamp 1698431365
transform 1 0 26544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A3
timestamp 1698431365
transform 1 0 31472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A4
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__B2
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__C2
timestamp 1698431365
transform -1 0 17920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A2
timestamp 1698431365
transform -1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A1
timestamp 1698431365
transform 1 0 23296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__S0
timestamp 1698431365
transform -1 0 26880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A1
timestamp 1698431365
transform -1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__A1
timestamp 1698431365
transform 1 0 39760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A2
timestamp 1698431365
transform 1 0 35056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__A2
timestamp 1698431365
transform 1 0 29344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A2
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1698431365
transform -1 0 6944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A1
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A2
timestamp 1698431365
transform 1 0 10640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A1
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A3
timestamp 1698431365
transform -1 0 10192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__B
timestamp 1698431365
transform -1 0 9408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1698431365
transform -1 0 16352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1698431365
transform -1 0 18928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A2
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A2
timestamp 1698431365
transform 1 0 40096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__I
timestamp 1698431365
transform 1 0 42000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A4
timestamp 1698431365
transform -1 0 41328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A2
timestamp 1698431365
transform 1 0 26992 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A2
timestamp 1698431365
transform 1 0 23744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__I
timestamp 1698431365
transform -1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1698431365
transform -1 0 26208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A2
timestamp 1698431365
transform 1 0 16240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A3
timestamp 1698431365
transform -1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__B2
timestamp 1698431365
transform -1 0 21504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__A1
timestamp 1698431365
transform 1 0 23744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__A1
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__B2
timestamp 1698431365
transform 1 0 32816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__A2
timestamp 1698431365
transform 1 0 37856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__B
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A2
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__B
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A1
timestamp 1698431365
transform -1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__A1
timestamp 1698431365
transform 1 0 38416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1958__A1
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__I
timestamp 1698431365
transform -1 0 22512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A2
timestamp 1698431365
transform -1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A2
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__B2
timestamp 1698431365
transform -1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__B
timestamp 1698431365
transform 1 0 43456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__I
timestamp 1698431365
transform -1 0 24416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A2
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A2
timestamp 1698431365
transform -1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__C
timestamp 1698431365
transform 1 0 28000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__A2
timestamp 1698431365
transform 1 0 29344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__B
timestamp 1698431365
transform -1 0 30016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__C
timestamp 1698431365
transform -1 0 32704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__A1
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__A2
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__B2
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A1
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A1
timestamp 1698431365
transform 1 0 32928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform -1 0 42112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__A2
timestamp 1698431365
transform -1 0 29120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A1
timestamp 1698431365
transform -1 0 30128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__B2
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__A1
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__A2
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__S
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A1
timestamp 1698431365
transform -1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__A1
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__A2
timestamp 1698431365
transform 1 0 19712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__B
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A2
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A1
timestamp 1698431365
transform -1 0 39088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A1
timestamp 1698431365
transform 1 0 43120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A2
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A1
timestamp 1698431365
transform 1 0 34832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__B
timestamp 1698431365
transform -1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__A2
timestamp 1698431365
transform -1 0 31136 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__A2
timestamp 1698431365
transform -1 0 31808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__C
timestamp 1698431365
transform 1 0 35392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__C
timestamp 1698431365
transform 1 0 47040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__A1
timestamp 1698431365
transform -1 0 36512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__A2
timestamp 1698431365
transform 1 0 36400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__B1
timestamp 1698431365
transform -1 0 37072 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__B2
timestamp 1698431365
transform 1 0 36176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__A2
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2105__A1
timestamp 1698431365
transform 1 0 33712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__A1
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A1
timestamp 1698431365
transform 1 0 43680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A1
timestamp 1698431365
transform 1 0 35728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__A1
timestamp 1698431365
transform 1 0 47376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A2
timestamp 1698431365
transform -1 0 17920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__I
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__A2
timestamp 1698431365
transform 1 0 18256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__I
timestamp 1698431365
transform -1 0 23520 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A2
timestamp 1698431365
transform 1 0 20272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__C
timestamp 1698431365
transform 1 0 19936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2199__I
timestamp 1698431365
transform 1 0 27888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A2
timestamp 1698431365
transform -1 0 21840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__A2
timestamp 1698431365
transform 1 0 28000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__A1
timestamp 1698431365
transform 1 0 26880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A1
timestamp 1698431365
transform 1 0 32592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__I
timestamp 1698431365
transform 1 0 14448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A2
timestamp 1698431365
transform 1 0 22736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A1
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A2
timestamp 1698431365
transform 1 0 31136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__B
timestamp 1698431365
transform 1 0 30688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__B
timestamp 1698431365
transform -1 0 14896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__A3
timestamp 1698431365
transform -1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__C
timestamp 1698431365
transform 1 0 19936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A2
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A2
timestamp 1698431365
transform -1 0 9296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__B2
timestamp 1698431365
transform -1 0 25536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A1
timestamp 1698431365
transform 1 0 25424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A1
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A2
timestamp 1698431365
transform -1 0 26880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__B1
timestamp 1698431365
transform 1 0 31696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__I
timestamp 1698431365
transform 1 0 29680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__B
timestamp 1698431365
transform 1 0 11200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__A2
timestamp 1698431365
transform 1 0 18368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__A1
timestamp 1698431365
transform 1 0 16800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A3
timestamp 1698431365
transform 1 0 19936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__A1
timestamp 1698431365
transform 1 0 16240 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__I
timestamp 1698431365
transform 1 0 27440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__A2
timestamp 1698431365
transform 1 0 25312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A2
timestamp 1698431365
transform 1 0 22064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__B
timestamp 1698431365
transform 1 0 38192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2273__A1
timestamp 1698431365
transform -1 0 41328 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__A1
timestamp 1698431365
transform -1 0 39872 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__A2
timestamp 1698431365
transform 1 0 20720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2277__A1
timestamp 1698431365
transform -1 0 21840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2277__B
timestamp 1698431365
transform -1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__B
timestamp 1698431365
transform -1 0 14672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A2
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1698431365
transform 1 0 35056 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__B
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__B
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A3
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__A1
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__A2
timestamp 1698431365
transform 1 0 30240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A1
timestamp 1698431365
transform -1 0 34720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A1
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__B
timestamp 1698431365
transform -1 0 11536 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A1
timestamp 1698431365
transform -1 0 28784 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A2
timestamp 1698431365
transform 1 0 29008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2324__A2
timestamp 1698431365
transform -1 0 19376 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__A3
timestamp 1698431365
transform -1 0 13888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__A2
timestamp 1698431365
transform 1 0 26544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__B2
timestamp 1698431365
transform -1 0 28224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A2
timestamp 1698431365
transform 1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__C
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1698431365
transform -1 0 22736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__B1
timestamp 1698431365
transform 1 0 20384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__A1
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__C1
timestamp 1698431365
transform 1 0 30688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A2
timestamp 1698431365
transform 1 0 39200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A2
timestamp 1698431365
transform -1 0 25424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A2
timestamp 1698431365
transform 1 0 16688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A2
timestamp 1698431365
transform 1 0 16352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A1
timestamp 1698431365
transform 1 0 15680 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__A2
timestamp 1698431365
transform -1 0 41552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A2
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2394__A2
timestamp 1698431365
transform 1 0 12320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A2
timestamp 1698431365
transform -1 0 16128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A2
timestamp 1698431365
transform 1 0 12320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A3
timestamp 1698431365
transform 1 0 14672 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__B
timestamp 1698431365
transform 1 0 15456 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__A2
timestamp 1698431365
transform 1 0 21504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__B
timestamp 1698431365
transform -1 0 13104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__B2
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__C
timestamp 1698431365
transform -1 0 10640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A1
timestamp 1698431365
transform -1 0 26768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__B1
timestamp 1698431365
transform 1 0 16240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2413__A2
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A2
timestamp 1698431365
transform -1 0 21056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A3
timestamp 1698431365
transform -1 0 21504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__A3
timestamp 1698431365
transform 1 0 23184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A2
timestamp 1698431365
transform 1 0 25312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__A2
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2433__A2
timestamp 1698431365
transform -1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A2
timestamp 1698431365
transform 1 0 26656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A4
timestamp 1698431365
transform 1 0 29232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1698431365
transform 1 0 28112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1698431365
transform 1 0 29680 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A2
timestamp 1698431365
transform -1 0 28112 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A2
timestamp 1698431365
transform -1 0 14448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A2
timestamp 1698431365
transform 1 0 38304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__B
timestamp 1698431365
transform 1 0 39648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__A2
timestamp 1698431365
transform 1 0 21392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__B1
timestamp 1698431365
transform 1 0 14560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__A2
timestamp 1698431365
transform 1 0 18368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2458__I
timestamp 1698431365
transform -1 0 16464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A2
timestamp 1698431365
transform 1 0 17360 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2460__A2
timestamp 1698431365
transform -1 0 20496 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A2
timestamp 1698431365
transform -1 0 37632 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__A1
timestamp 1698431365
transform -1 0 18592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A2
timestamp 1698431365
transform 1 0 26096 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A3
timestamp 1698431365
transform 1 0 25648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__S
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2494__A2
timestamp 1698431365
transform 1 0 15568 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A2
timestamp 1698431365
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A2
timestamp 1698431365
transform -1 0 11760 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A3
timestamp 1698431365
transform -1 0 11312 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1698431365
transform 1 0 12880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A2
timestamp 1698431365
transform -1 0 14784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__I0
timestamp 1698431365
transform 1 0 40432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A4
timestamp 1698431365
transform 1 0 33824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__A2
timestamp 1698431365
transform 1 0 22288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__A2
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A2
timestamp 1698431365
transform -1 0 22176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__B2
timestamp 1698431365
transform 1 0 21504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A2
timestamp 1698431365
transform -1 0 30464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2523__B
timestamp 1698431365
transform 1 0 35168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__A2
timestamp 1698431365
transform -1 0 40208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__B
timestamp 1698431365
transform -1 0 37856 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A1
timestamp 1698431365
transform -1 0 14672 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A2
timestamp 1698431365
transform 1 0 15680 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A1
timestamp 1698431365
transform 1 0 16912 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A2
timestamp 1698431365
transform -1 0 15568 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__B
timestamp 1698431365
transform 1 0 17472 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A2
timestamp 1698431365
transform 1 0 20160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__A1
timestamp 1698431365
transform -1 0 24192 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A2
timestamp 1698431365
transform -1 0 39088 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__I
timestamp 1698431365
transform -1 0 33488 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__I
timestamp 1698431365
transform -1 0 16576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__A3
timestamp 1698431365
transform -1 0 16128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A1
timestamp 1698431365
transform 1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A2
timestamp 1698431365
transform -1 0 19264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A2
timestamp 1698431365
transform -1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__B1
timestamp 1698431365
transform 1 0 23296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__A2
timestamp 1698431365
transform 1 0 26432 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__A1
timestamp 1698431365
transform 1 0 26432 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__B
timestamp 1698431365
transform 1 0 28112 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__C
timestamp 1698431365
transform 1 0 29232 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__A3
timestamp 1698431365
transform 1 0 20720 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A2
timestamp 1698431365
transform 1 0 24528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__C
timestamp 1698431365
transform -1 0 26544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__A1
timestamp 1698431365
transform -1 0 39984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__A2
timestamp 1698431365
transform 1 0 23520 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__A1
timestamp 1698431365
transform 1 0 19488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__A3
timestamp 1698431365
transform 1 0 19040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__A1
timestamp 1698431365
transform 1 0 21168 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__I
timestamp 1698431365
transform 1 0 40992 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__A1
timestamp 1698431365
transform 1 0 21392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__A3
timestamp 1698431365
transform -1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__A4
timestamp 1698431365
transform -1 0 22288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A1
timestamp 1698431365
transform 1 0 15680 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__B
timestamp 1698431365
transform 1 0 17472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__B
timestamp 1698431365
transform -1 0 18704 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A2
timestamp 1698431365
transform -1 0 18480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__B1
timestamp 1698431365
transform 1 0 18704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A1
timestamp 1698431365
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A2
timestamp 1698431365
transform 1 0 32144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__A2
timestamp 1698431365
transform -1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A1
timestamp 1698431365
transform -1 0 18816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A2
timestamp 1698431365
transform -1 0 19264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A1
timestamp 1698431365
transform 1 0 25760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__A1
timestamp 1698431365
transform 1 0 26880 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__A2
timestamp 1698431365
transform -1 0 31136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__A1
timestamp 1698431365
transform -1 0 27776 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__A2
timestamp 1698431365
transform 1 0 28784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__A1
timestamp 1698431365
transform 1 0 29232 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A2
timestamp 1698431365
transform 1 0 27440 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__A1
timestamp 1698431365
transform 1 0 28560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__C
timestamp 1698431365
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__A2
timestamp 1698431365
transform -1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__B2
timestamp 1698431365
transform 1 0 29232 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__A1
timestamp 1698431365
transform 1 0 30464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__A2
timestamp 1698431365
transform 1 0 43904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__A1
timestamp 1698431365
transform -1 0 45136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A1
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A2
timestamp 1698431365
transform -1 0 25760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__A1
timestamp 1698431365
transform -1 0 11872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__A1
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__A1
timestamp 1698431365
transform 1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A1
timestamp 1698431365
transform 1 0 20272 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__A1
timestamp 1698431365
transform 1 0 18816 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__A1
timestamp 1698431365
transform -1 0 24528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__A1
timestamp 1698431365
transform -1 0 24752 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2748__A1
timestamp 1698431365
transform -1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__A1
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__A2
timestamp 1698431365
transform -1 0 23520 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2750__A1
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__A1
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__A1
timestamp 1698431365
transform 1 0 26432 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2758__A1
timestamp 1698431365
transform -1 0 19264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A1
timestamp 1698431365
transform 1 0 21392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A1
timestamp 1698431365
transform -1 0 27552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A2
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2768__A2
timestamp 1698431365
transform -1 0 22960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2772__A1
timestamp 1698431365
transform 1 0 23744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__D
timestamp 1698431365
transform 1 0 45360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2782__D
timestamp 1698431365
transform -1 0 35728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2787__CLK
timestamp 1698431365
transform -1 0 19040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__CLK
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout44_I
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout53_I
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout58_I
timestamp 1698431365
transform 1 0 10304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout64_I
timestamp 1698431365
transform 1 0 27888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout68_I
timestamp 1698431365
transform 1 0 5712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout69_I
timestamp 1698431365
transform 1 0 4368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout70_I
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 57680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1698431365
transform -1 0 4928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout44
timestamp 1698431365
transform -1 0 33600 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout45
timestamp 1698431365
transform -1 0 32368 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout46
timestamp 1698431365
transform -1 0 41552 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout47
timestamp 1698431365
transform -1 0 42448 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout48
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout49
timestamp 1698431365
transform 1 0 33040 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout50
timestamp 1698431365
transform -1 0 33936 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout51
timestamp 1698431365
transform -1 0 18144 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout52
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout53
timestamp 1698431365
transform -1 0 31248 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout54
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout55
timestamp 1698431365
transform 1 0 10192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout56
timestamp 1698431365
transform -1 0 10080 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout57
timestamp 1698431365
transform 1 0 9408 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout58
timestamp 1698431365
transform 1 0 8736 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout59
timestamp 1698431365
transform -1 0 28784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout60
timestamp 1698431365
transform -1 0 37408 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout61
timestamp 1698431365
transform -1 0 41776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout62
timestamp 1698431365
transform -1 0 45360 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout63
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout64
timestamp 1698431365
transform 1 0 28112 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout65
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1698431365
transform 1 0 3920 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout67
timestamp 1698431365
transform -1 0 6496 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout68
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout69
timestamp 1698431365
transform 1 0 4592 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout70
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_41
timestamp 1698431365
transform 1 0 5936 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_53 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_59
timestamp 1698431365
transform 1 0 7952 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_78
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_82
timestamp 1698431365
transform 1 0 10528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_86
timestamp 1698431365
transform 1 0 10976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_90
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_94
timestamp 1698431365
transform 1 0 11872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_98
timestamp 1698431365
transform 1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_112
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_116
timestamp 1698431365
transform 1 0 14336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_120
timestamp 1698431365
transform 1 0 14784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_124
timestamp 1698431365
transform 1 0 15232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_128
timestamp 1698431365
transform 1 0 15680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_132
timestamp 1698431365
transform 1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_148
timestamp 1698431365
transform 1 0 17920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_154
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_158
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_162
timestamp 1698431365
transform 1 0 19488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_166
timestamp 1698431365
transform 1 0 19936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_176
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_179
timestamp 1698431365
transform 1 0 21392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_191
timestamp 1698431365
transform 1 0 22736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_214
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_216
timestamp 1698431365
transform 1 0 25536 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_229
timestamp 1698431365
transform 1 0 26992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_233
timestamp 1698431365
transform 1 0 27440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_248
timestamp 1698431365
transform 1 0 29120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_260
timestamp 1698431365
transform 1 0 30464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_264
timestamp 1698431365
transform 1 0 30912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_268
timestamp 1698431365
transform 1 0 31360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_278
timestamp 1698431365
transform 1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_282
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_286
timestamp 1698431365
transform 1 0 33376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_290
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_294
timestamp 1698431365
transform 1 0 34272 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_302
timestamp 1698431365
transform 1 0 35168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_414
timestamp 1698431365
transform 1 0 47712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_448
timestamp 1698431365
transform 1 0 51520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_498
timestamp 1698431365
transform 1 0 57120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_500
timestamp 1698431365
transform 1 0 57344 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_74
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_77
timestamp 1698431365
transform 1 0 9968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_81
timestamp 1698431365
transform 1 0 10416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_85
timestamp 1698431365
transform 1 0 10864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_89
timestamp 1698431365
transform 1 0 11312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_99
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_117
timestamp 1698431365
transform 1 0 14448 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_126
timestamp 1698431365
transform 1 0 15456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_152
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_163
timestamp 1698431365
transform 1 0 19600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_238
timestamp 1698431365
transform 1 0 28000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_258
timestamp 1698431365
transform 1 0 30240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_273
timestamp 1698431365
transform 1 0 31920 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_290
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_294
timestamp 1698431365
transform 1 0 34272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_298
timestamp 1698431365
transform 1 0 34720 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_330
timestamp 1698431365
transform 1 0 38304 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_358
timestamp 1698431365
transform 1 0 41440 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_390
timestamp 1698431365
transform 1 0 45024 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_398
timestamp 1698431365
transform 1 0 45920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_418
timestamp 1698431365
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_500
timestamp 1698431365
transform 1 0 57344 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_504
timestamp 1698431365
transform 1 0 57792 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_71
timestamp 1698431365
transform 1 0 9296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_75
timestamp 1698431365
transform 1 0 9744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_85
timestamp 1698431365
transform 1 0 10864 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_94
timestamp 1698431365
transform 1 0 11872 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_117
timestamp 1698431365
transform 1 0 14448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_129
timestamp 1698431365
transform 1 0 15792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_131
timestamp 1698431365
transform 1 0 16016 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_146
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_156
timestamp 1698431365
transform 1 0 18816 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_186
timestamp 1698431365
transform 1 0 22176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_215
timestamp 1698431365
transform 1 0 25424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_217
timestamp 1698431365
transform 1 0 25648 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_228
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_283
timestamp 1698431365
transform 1 0 33040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_287
timestamp 1698431365
transform 1 0 33488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_291
timestamp 1698431365
transform 1 0 33936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_295
timestamp 1698431365
transform 1 0 34384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_299
timestamp 1698431365
transform 1 0 34832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_302
timestamp 1698431365
transform 1 0 35168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_306
timestamp 1698431365
transform 1 0 35616 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_358
timestamp 1698431365
transform 1 0 41440 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_389
timestamp 1698431365
transform 1 0 44912 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_425
timestamp 1698431365
transform 1 0 48944 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_441
timestamp 1698431365
transform 1 0 50736 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_449
timestamp 1698431365
transform 1 0 51632 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_453
timestamp 1698431365
transform 1 0 52080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_34
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_50
timestamp 1698431365
transform 1 0 6944 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_54
timestamp 1698431365
transform 1 0 7392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_58
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 9632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_85
timestamp 1698431365
transform 1 0 10864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_87
timestamp 1698431365
transform 1 0 11088 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_90
timestamp 1698431365
transform 1 0 11424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_94
timestamp 1698431365
transform 1 0 11872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_126
timestamp 1698431365
transform 1 0 15456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_132
timestamp 1698431365
transform 1 0 16128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_151
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_162
timestamp 1698431365
transform 1 0 19488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_242
timestamp 1698431365
transform 1 0 28448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_307
timestamp 1698431365
transform 1 0 35728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_311
timestamp 1698431365
transform 1 0 36176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_315
timestamp 1698431365
transform 1 0 36624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_319
timestamp 1698431365
transform 1 0 37072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_323
timestamp 1698431365
transform 1 0 37520 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_356
timestamp 1698431365
transform 1 0 41216 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_370
timestamp 1698431365
transform 1 0 42784 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_413
timestamp 1698431365
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_417
timestamp 1698431365
transform 1 0 48048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_500
timestamp 1698431365
transform 1 0 57344 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_504
timestamp 1698431365
transform 1 0 57792 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_49
timestamp 1698431365
transform 1 0 6832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_51
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_54
timestamp 1698431365
transform 1 0 7392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_66
timestamp 1698431365
transform 1 0 8736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_122
timestamp 1698431365
transform 1 0 15008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_140
timestamp 1698431365
transform 1 0 17024 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_238
timestamp 1698431365
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_257
timestamp 1698431365
transform 1 0 30128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_259
timestamp 1698431365
transform 1 0 30352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_300
timestamp 1698431365
transform 1 0 34944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_304
timestamp 1698431365
transform 1 0 35392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_308
timestamp 1698431365
transform 1 0 35840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_312
timestamp 1698431365
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_329
timestamp 1698431365
transform 1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_333
timestamp 1698431365
transform 1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_335
timestamp 1698431365
transform 1 0 38864 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_338
timestamp 1698431365
transform 1 0 39200 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_346
timestamp 1698431365
transform 1 0 40096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_373
timestamp 1698431365
transform 1 0 43120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_377
timestamp 1698431365
transform 1 0 43568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_400
timestamp 1698431365
transform 1 0 46144 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_408
timestamp 1698431365
transform 1 0 47040 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_435
timestamp 1698431365
transform 1 0 50064 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_454
timestamp 1698431365
transform 1 0 52192 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_42
timestamp 1698431365
transform 1 0 6048 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_46
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_54
timestamp 1698431365
transform 1 0 7392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_82
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_103
timestamp 1698431365
transform 1 0 12880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_137
timestamp 1698431365
transform 1 0 16688 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_149
timestamp 1698431365
transform 1 0 18032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_151
timestamp 1698431365
transform 1 0 18256 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_160
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_166
timestamp 1698431365
transform 1 0 19936 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_175
timestamp 1698431365
transform 1 0 20944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_177
timestamp 1698431365
transform 1 0 21168 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_180
timestamp 1698431365
transform 1 0 21504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_225
timestamp 1698431365
transform 1 0 26544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_254
timestamp 1698431365
transform 1 0 29792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_299
timestamp 1698431365
transform 1 0 34832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_335
timestamp 1698431365
transform 1 0 38864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_337
timestamp 1698431365
transform 1 0 39088 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_344
timestamp 1698431365
transform 1 0 39872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_348
timestamp 1698431365
transform 1 0 40320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_365
timestamp 1698431365
transform 1 0 42224 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_373
timestamp 1698431365
transform 1 0 43120 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_401
timestamp 1698431365
transform 1 0 46256 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_417
timestamp 1698431365
transform 1 0 48048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_419
timestamp 1698431365
transform 1 0 48272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_430
timestamp 1698431365
transform 1 0 49504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_451
timestamp 1698431365
transform 1 0 51856 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_483
timestamp 1698431365
transform 1 0 55440 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_487
timestamp 1698431365
transform 1 0 55888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_489
timestamp 1698431365
transform 1 0 56112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_58
timestamp 1698431365
transform 1 0 7840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_74
timestamp 1698431365
transform 1 0 9632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_78
timestamp 1698431365
transform 1 0 10080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_225
timestamp 1698431365
transform 1 0 26544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_249
timestamp 1698431365
transform 1 0 29232 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_252
timestamp 1698431365
transform 1 0 29568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_256
timestamp 1698431365
transform 1 0 30016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_298
timestamp 1698431365
transform 1 0 34720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_302
timestamp 1698431365
transform 1 0 35168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_310
timestamp 1698431365
transform 1 0 36064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_333
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_341
timestamp 1698431365
transform 1 0 39536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_345
timestamp 1698431365
transform 1 0 39984 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_358
timestamp 1698431365
transform 1 0 41440 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_374
timestamp 1698431365
transform 1 0 43232 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_382
timestamp 1698431365
transform 1 0 44128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_403
timestamp 1698431365
transform 1 0 46480 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_411
timestamp 1698431365
transform 1 0 47376 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_430
timestamp 1698431365
transform 1 0 49504 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_446
timestamp 1698431365
transform 1 0 51296 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_473
timestamp 1698431365
transform 1 0 54320 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_481
timestamp 1698431365
transform 1 0 55216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_6
timestamp 1698431365
transform 1 0 2016 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_38
timestamp 1698431365
transform 1 0 5600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_44
timestamp 1698431365
transform 1 0 6272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_65
timestamp 1698431365
transform 1 0 8624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_125
timestamp 1698431365
transform 1 0 15344 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_165
timestamp 1698431365
transform 1 0 19824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_169
timestamp 1698431365
transform 1 0 20272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_187
timestamp 1698431365
transform 1 0 22288 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_295
timestamp 1698431365
transform 1 0 34384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_299
timestamp 1698431365
transform 1 0 34832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_339
timestamp 1698431365
transform 1 0 39312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_343
timestamp 1698431365
transform 1 0 39760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_345
timestamp 1698431365
transform 1 0 39984 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_365
timestamp 1698431365
transform 1 0 42224 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_371
timestamp 1698431365
transform 1 0 42896 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_391
timestamp 1698431365
transform 1 0 45136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_397
timestamp 1698431365
transform 1 0 45808 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_413
timestamp 1698431365
transform 1 0 47600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_417
timestamp 1698431365
transform 1 0 48048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_427
timestamp 1698431365
transform 1 0 49168 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_443
timestamp 1698431365
transform 1 0 50960 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_451
timestamp 1698431365
transform 1 0 51856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_453
timestamp 1698431365
transform 1 0 52080 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_472
timestamp 1698431365
transform 1 0 54208 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_488
timestamp 1698431365
transform 1 0 56000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_39
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_42
timestamp 1698431365
transform 1 0 6048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_46
timestamp 1698431365
transform 1 0 6496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_50
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_95
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_197
timestamp 1698431365
transform 1 0 23408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_199
timestamp 1698431365
transform 1 0 23632 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_210
timestamp 1698431365
transform 1 0 24864 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_249
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_301
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_305
timestamp 1698431365
transform 1 0 35504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_333
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_337
timestamp 1698431365
transform 1 0 39088 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_374
timestamp 1698431365
transform 1 0 43232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_399
timestamp 1698431365
transform 1 0 46032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_413
timestamp 1698431365
transform 1 0 47600 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_427
timestamp 1698431365
transform 1 0 49168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_435
timestamp 1698431365
transform 1 0 50064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_437
timestamp 1698431365
transform 1 0 50288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_453
timestamp 1698431365
transform 1 0 52080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_36
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_76
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_199
timestamp 1698431365
transform 1 0 23632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_230
timestamp 1698431365
transform 1 0 27104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_232
timestamp 1698431365
transform 1 0 27328 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_264
timestamp 1698431365
transform 1 0 30912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_266
timestamp 1698431365
transform 1 0 31136 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_299
timestamp 1698431365
transform 1 0 34832 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_303
timestamp 1698431365
transform 1 0 35280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_342
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_358
timestamp 1698431365
transform 1 0 41440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_362
timestamp 1698431365
transform 1 0 41888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_366
timestamp 1698431365
transform 1 0 42336 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_378
timestamp 1698431365
transform 1 0 43680 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_386
timestamp 1698431365
transform 1 0 44576 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_430
timestamp 1698431365
transform 1 0 49504 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_453
timestamp 1698431365
transform 1 0 52080 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_457
timestamp 1698431365
transform 1 0 52528 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_464
timestamp 1698431365
transform 1 0 53312 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_471
timestamp 1698431365
transform 1 0 54096 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_487
timestamp 1698431365
transform 1 0 55888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_489
timestamp 1698431365
transform 1 0 56112 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_48
timestamp 1698431365
transform 1 0 6720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_52
timestamp 1698431365
transform 1 0 7168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_56
timestamp 1698431365
transform 1 0 7616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_60
timestamp 1698431365
transform 1 0 8064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_64
timestamp 1698431365
transform 1 0 8512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_68
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_72
timestamp 1698431365
transform 1 0 9408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_76
timestamp 1698431365
transform 1 0 9856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_80
timestamp 1698431365
transform 1 0 10304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_152
timestamp 1698431365
transform 1 0 18368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_154
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_257
timestamp 1698431365
transform 1 0 30128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_265
timestamp 1698431365
transform 1 0 31024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_337
timestamp 1698431365
transform 1 0 39088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_341
timestamp 1698431365
transform 1 0 39536 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_345
timestamp 1698431365
transform 1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_349
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_353
timestamp 1698431365
transform 1 0 40880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_357
timestamp 1698431365
transform 1 0 41328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_399
timestamp 1698431365
transform 1 0 46032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_401
timestamp 1698431365
transform 1 0 46256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_422
timestamp 1698431365
transform 1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_424
timestamp 1698431365
transform 1 0 48832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_435
timestamp 1698431365
transform 1 0 50064 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_476
timestamp 1698431365
transform 1 0 54656 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_508
timestamp 1698431365
transform 1 0 58240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_46
timestamp 1698431365
transform 1 0 6496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_65
timestamp 1698431365
transform 1 0 8624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_74
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_131
timestamp 1698431365
transform 1 0 16016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_308
timestamp 1698431365
transform 1 0 35840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_328
timestamp 1698431365
transform 1 0 38080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_332
timestamp 1698431365
transform 1 0 38528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_334
timestamp 1698431365
transform 1 0 38752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_343
timestamp 1698431365
transform 1 0 39760 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_354
timestamp 1698431365
transform 1 0 40992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_402
timestamp 1698431365
transform 1 0 46368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_404
timestamp 1698431365
transform 1 0 46592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_448
timestamp 1698431365
transform 1 0 51520 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_468
timestamp 1698431365
transform 1 0 53760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_470
timestamp 1698431365
transform 1 0 53984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_489
timestamp 1698431365
transform 1 0 56112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_109
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_118
timestamp 1698431365
transform 1 0 14560 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_215
timestamp 1698431365
transform 1 0 25424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_217
timestamp 1698431365
transform 1 0 25648 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_298
timestamp 1698431365
transform 1 0 34720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_302
timestamp 1698431365
transform 1 0 35168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_364
timestamp 1698431365
transform 1 0 42112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_368
timestamp 1698431365
transform 1 0 42560 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_395
timestamp 1698431365
transform 1 0 45584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_399
timestamp 1698431365
transform 1 0 46032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_401
timestamp 1698431365
transform 1 0 46256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_410
timestamp 1698431365
transform 1 0 47264 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_426
timestamp 1698431365
transform 1 0 49056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_434
timestamp 1698431365
transform 1 0 49952 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_469
timestamp 1698431365
transform 1 0 53872 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_477
timestamp 1698431365
transform 1 0 54768 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_481
timestamp 1698431365
transform 1 0 55216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_38
timestamp 1698431365
transform 1 0 5600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_48
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_115
timestamp 1698431365
transform 1 0 14224 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_154
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_190
timestamp 1698431365
transform 1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_221
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_256
timestamp 1698431365
transform 1 0 30016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_356
timestamp 1698431365
transform 1 0 41216 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_380
timestamp 1698431365
transform 1 0 43904 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_388
timestamp 1698431365
transform 1 0 44800 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_401
timestamp 1698431365
transform 1 0 46256 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_438
timestamp 1698431365
transform 1 0 50400 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_446
timestamp 1698431365
transform 1 0 51296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_448
timestamp 1698431365
transform 1 0 51520 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_456
timestamp 1698431365
transform 1 0 52416 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_488
timestamp 1698431365
transform 1 0 56000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_41
timestamp 1698431365
transform 1 0 5936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_69
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_195
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_302
timestamp 1698431365
transform 1 0 35168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_308
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_379
timestamp 1698431365
transform 1 0 43792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_418
timestamp 1698431365
transform 1 0 48160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_444
timestamp 1698431365
transform 1 0 51072 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_452
timestamp 1698431365
transform 1 0 51968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_454
timestamp 1698431365
transform 1 0 52192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_465
timestamp 1698431365
transform 1 0 53424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_469
timestamp 1698431365
transform 1 0 53872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_477
timestamp 1698431365
transform 1 0 54768 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_481
timestamp 1698431365
transform 1 0 55216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_36
timestamp 1698431365
transform 1 0 5376 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_39
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_126
timestamp 1698431365
transform 1 0 15456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_128
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_161
timestamp 1698431365
transform 1 0 19376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_242
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_244
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_292
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_302
timestamp 1698431365
transform 1 0 35168 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_306
timestamp 1698431365
transform 1 0 35616 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_322
timestamp 1698431365
transform 1 0 37408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_341
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_354
timestamp 1698431365
transform 1 0 40992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_357
timestamp 1698431365
transform 1 0 41328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_361
timestamp 1698431365
transform 1 0 41776 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_377
timestamp 1698431365
transform 1 0 43568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_393
timestamp 1698431365
transform 1 0 45360 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_397
timestamp 1698431365
transform 1 0 45808 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_400
timestamp 1698431365
transform 1 0 46144 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_447
timestamp 1698431365
transform 1 0 51408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_455
timestamp 1698431365
transform 1 0 52304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_474
timestamp 1698431365
transform 1 0 54432 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_47
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_53
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_73
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_86
timestamp 1698431365
transform 1 0 10976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_90
timestamp 1698431365
transform 1 0 11424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_97
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_279
timestamp 1698431365
transform 1 0 32592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_281
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_371
timestamp 1698431365
transform 1 0 42896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_375
timestamp 1698431365
transform 1 0 43344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_377
timestamp 1698431365
transform 1 0 43568 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_393
timestamp 1698431365
transform 1 0 45360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_397
timestamp 1698431365
transform 1 0 45808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_420
timestamp 1698431365
transform 1 0 48384 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_428
timestamp 1698431365
transform 1 0 49280 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_433
timestamp 1698431365
transform 1 0 49840 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_441
timestamp 1698431365
transform 1 0 50736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_445
timestamp 1698431365
transform 1 0 51184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_470
timestamp 1698431365
transform 1 0 53984 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_502
timestamp 1698431365
transform 1 0 57568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_506
timestamp 1698431365
transform 1 0 58016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_508
timestamp 1698431365
transform 1 0 58240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_26
timestamp 1698431365
transform 1 0 4256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_59
timestamp 1698431365
transform 1 0 7952 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_61
timestamp 1698431365
transform 1 0 8176 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_275
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_297
timestamp 1698431365
transform 1 0 34608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_304
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_312
timestamp 1698431365
transform 1 0 36288 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_316
timestamp 1698431365
transform 1 0 36736 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_325
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_345
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_365
timestamp 1698431365
transform 1 0 42224 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_381
timestamp 1698431365
transform 1 0 44016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_410
timestamp 1698431365
transform 1 0 47264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_418
timestamp 1698431365
transform 1 0 48160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_454
timestamp 1698431365
transform 1 0 52192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_458
timestamp 1698431365
transform 1 0 52640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_460
timestamp 1698431365
transform 1 0 52864 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_483
timestamp 1698431365
transform 1 0 55440 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_487
timestamp 1698431365
transform 1 0 55888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_489
timestamp 1698431365
transform 1 0 56112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_6
timestamp 1698431365
transform 1 0 2016 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_22
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_57
timestamp 1698431365
transform 1 0 7728 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_60
timestamp 1698431365
transform 1 0 8064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_64
timestamp 1698431365
transform 1 0 8512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_68
timestamp 1698431365
transform 1 0 8960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_80
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_84
timestamp 1698431365
transform 1 0 10752 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_96
timestamp 1698431365
transform 1 0 12096 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_131
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_190
timestamp 1698431365
transform 1 0 22624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_192
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_195
timestamp 1698431365
transform 1 0 23184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_216
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_220
timestamp 1698431365
transform 1 0 25984 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_223
timestamp 1698431365
transform 1 0 26320 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_227
timestamp 1698431365
transform 1 0 26768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_231
timestamp 1698431365
transform 1 0 27216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_235
timestamp 1698431365
transform 1 0 27664 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_267
timestamp 1698431365
transform 1 0 31248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_271
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_280
timestamp 1698431365
transform 1 0 32704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_302
timestamp 1698431365
transform 1 0 35168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_308
timestamp 1698431365
transform 1 0 35840 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_327
timestamp 1698431365
transform 1 0 37968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_344
timestamp 1698431365
transform 1 0 39872 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_348
timestamp 1698431365
transform 1 0 40320 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_350
timestamp 1698431365
transform 1 0 40544 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_372
timestamp 1698431365
transform 1 0 43008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_380
timestamp 1698431365
transform 1 0 43904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_389
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_396
timestamp 1698431365
transform 1 0 45696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_400
timestamp 1698431365
transform 1 0 46144 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_415
timestamp 1698431365
transform 1 0 47824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_423
timestamp 1698431365
transform 1 0 48720 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_432
timestamp 1698431365
transform 1 0 49728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_446
timestamp 1698431365
transform 1 0 51296 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698431365
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_482
timestamp 1698431365
transform 1 0 55328 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_42
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_46
timestamp 1698431365
transform 1 0 6496 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_61
timestamp 1698431365
transform 1 0 8176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_152
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_197
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_224
timestamp 1698431365
transform 1 0 26432 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_267
timestamp 1698431365
transform 1 0 31248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_271
timestamp 1698431365
transform 1 0 31696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_293
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_299
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_305
timestamp 1698431365
transform 1 0 35504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_309
timestamp 1698431365
transform 1 0 35952 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_325
timestamp 1698431365
transform 1 0 37744 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_390
timestamp 1698431365
transform 1 0 45024 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_415
timestamp 1698431365
transform 1 0 47824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_435
timestamp 1698431365
transform 1 0 50064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_437
timestamp 1698431365
transform 1 0 50288 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_6
timestamp 1698431365
transform 1 0 2016 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_22
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_57
timestamp 1698431365
transform 1 0 7728 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_63
timestamp 1698431365
transform 1 0 8400 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_99
timestamp 1698431365
transform 1 0 12432 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_151
timestamp 1698431365
transform 1 0 18256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_221
timestamp 1698431365
transform 1 0 26096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_266
timestamp 1698431365
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_268
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_302
timestamp 1698431365
transform 1 0 35168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_306
timestamp 1698431365
transform 1 0 35616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_349
timestamp 1698431365
transform 1 0 40432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_357
timestamp 1698431365
transform 1 0 41328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_364
timestamp 1698431365
transform 1 0 42112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_380
timestamp 1698431365
transform 1 0 43904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_397
timestamp 1698431365
transform 1 0 45808 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_414
timestamp 1698431365
transform 1 0 47712 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_430
timestamp 1698431365
transform 1 0 49504 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_434
timestamp 1698431365
transform 1 0 49952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_436
timestamp 1698431365
transform 1 0 50176 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_453
timestamp 1698431365
transform 1 0 52080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_470
timestamp 1698431365
transform 1 0 53984 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_502
timestamp 1698431365
transform 1 0 57568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_506
timestamp 1698431365
transform 1 0 58016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_508
timestamp 1698431365
transform 1 0 58240 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_34
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_48
timestamp 1698431365
transform 1 0 6720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_120
timestamp 1698431365
transform 1 0 14784 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_130
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_132
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_240
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_244
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_274
timestamp 1698431365
transform 1 0 32032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_294
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_331
timestamp 1698431365
transform 1 0 38416 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_358
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_367
timestamp 1698431365
transform 1 0 42448 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_399
timestamp 1698431365
transform 1 0 46032 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_415
timestamp 1698431365
transform 1 0 47824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_62
timestamp 1698431365
transform 1 0 8288 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_78
timestamp 1698431365
transform 1 0 10080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_82
timestamp 1698431365
transform 1 0 10528 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_85
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_89
timestamp 1698431365
transform 1 0 11312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_93
timestamp 1698431365
transform 1 0 11760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_151
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_190
timestamp 1698431365
transform 1 0 22624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_194
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_198
timestamp 1698431365
transform 1 0 23520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_202
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_204
timestamp 1698431365
transform 1 0 24192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_218
timestamp 1698431365
transform 1 0 25760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_222
timestamp 1698431365
transform 1 0 26208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_224
timestamp 1698431365
transform 1 0 26432 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_227
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_249
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_252
timestamp 1698431365
transform 1 0 29568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_261
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_274
timestamp 1698431365
transform 1 0 32032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_278
timestamp 1698431365
transform 1 0 32480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_280
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_333
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_352
timestamp 1698431365
transform 1 0 40768 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_356
timestamp 1698431365
transform 1 0 41216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_371
timestamp 1698431365
transform 1 0 42896 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_399
timestamp 1698431365
transform 1 0 46032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_416
timestamp 1698431365
transform 1 0 47936 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_424
timestamp 1698431365
transform 1 0 48832 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_452
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_461
timestamp 1698431365
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_463
timestamp 1698431365
transform 1 0 53200 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_482
timestamp 1698431365
transform 1 0 55328 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_28
timestamp 1698431365
transform 1 0 4480 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_36
timestamp 1698431365
transform 1 0 5376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_52
timestamp 1698431365
transform 1 0 7168 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_86
timestamp 1698431365
transform 1 0 10976 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_108
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698431365
transform 1 0 16240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_176
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_228
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_230
timestamp 1698431365
transform 1 0 27104 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_236
timestamp 1698431365
transform 1 0 27776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_273
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_301
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_305
timestamp 1698431365
transform 1 0 35504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_334
timestamp 1698431365
transform 1 0 38752 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_374
timestamp 1698431365
transform 1 0 43232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_390
timestamp 1698431365
transform 1 0 45024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_398
timestamp 1698431365
transform 1 0 45920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_402
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_424
timestamp 1698431365
transform 1 0 48832 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_454
timestamp 1698431365
transform 1 0 52192 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_458
timestamp 1698431365
transform 1 0 52640 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_478
timestamp 1698431365
transform 1 0 54880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_53
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_61
timestamp 1698431365
transform 1 0 8176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_98
timestamp 1698431365
transform 1 0 12320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_102
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_154
timestamp 1698431365
transform 1 0 18592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_156
timestamp 1698431365
transform 1 0 18816 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_223
timestamp 1698431365
transform 1 0 26320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_227
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_251
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_253
timestamp 1698431365
transform 1 0 29680 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_273
timestamp 1698431365
transform 1 0 31920 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_277
timestamp 1698431365
transform 1 0 32368 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_298
timestamp 1698431365
transform 1 0 34720 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_307
timestamp 1698431365
transform 1 0 35728 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_323
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_330
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_334
timestamp 1698431365
transform 1 0 38752 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_349
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_353
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_366
timestamp 1698431365
transform 1 0 42336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_370
timestamp 1698431365
transform 1 0 42784 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_402
timestamp 1698431365
transform 1 0 46368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_419
timestamp 1698431365
transform 1 0 48272 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_443
timestamp 1698431365
transform 1 0 50960 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_477
timestamp 1698431365
transform 1 0 54768 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_28
timestamp 1698431365
transform 1 0 4480 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_48
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_102
timestamp 1698431365
transform 1 0 12768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_160
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_181
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_189
timestamp 1698431365
transform 1 0 22512 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_204
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_219
timestamp 1698431365
transform 1 0 25872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_230
timestamp 1698431365
transform 1 0 27104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_263
timestamp 1698431365
transform 1 0 30800 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_272
timestamp 1698431365
transform 1 0 31808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_288
timestamp 1698431365
transform 1 0 33600 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_300
timestamp 1698431365
transform 1 0 34944 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_306
timestamp 1698431365
transform 1 0 35616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_310
timestamp 1698431365
transform 1 0 36064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_313
timestamp 1698431365
transform 1 0 36400 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_347
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_371
timestamp 1698431365
transform 1 0 42896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_375
timestamp 1698431365
transform 1 0 43344 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_400
timestamp 1698431365
transform 1 0 46144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_408
timestamp 1698431365
transform 1 0 47040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_410
timestamp 1698431365
transform 1 0 47264 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_413
timestamp 1698431365
transform 1 0 47600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_417
timestamp 1698431365
transform 1 0 48048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_431
timestamp 1698431365
transform 1 0 49616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_439
timestamp 1698431365
transform 1 0 50512 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_476
timestamp 1698431365
transform 1 0 54656 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_484
timestamp 1698431365
transform 1 0 55552 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_488
timestamp 1698431365
transform 1 0 56000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_59
timestamp 1698431365
transform 1 0 7952 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_67
timestamp 1698431365
transform 1 0 8848 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_76
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_80
timestamp 1698431365
transform 1 0 10304 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_91
timestamp 1698431365
transform 1 0 11536 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_109
timestamp 1698431365
transform 1 0 13552 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_118
timestamp 1698431365
transform 1 0 14560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_202
timestamp 1698431365
transform 1 0 23968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_206
timestamp 1698431365
transform 1 0 24416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_218
timestamp 1698431365
transform 1 0 25760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_266
timestamp 1698431365
transform 1 0 31136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_357
timestamp 1698431365
transform 1 0 41328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_361
timestamp 1698431365
transform 1 0 41776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_378
timestamp 1698431365
transform 1 0 43680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_411
timestamp 1698431365
transform 1 0 47376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_438
timestamp 1698431365
transform 1 0 50400 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_454
timestamp 1698431365
transform 1 0 52192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_479
timestamp 1698431365
transform 1 0 54992 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_30
timestamp 1698431365
transform 1 0 4704 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698431365
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_96
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_102
timestamp 1698431365
transform 1 0 12768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_110
timestamp 1698431365
transform 1 0 13664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698431365
transform 1 0 18144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_152
timestamp 1698431365
transform 1 0 18368 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_155
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_159
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_163
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_172
timestamp 1698431365
transform 1 0 20608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_176
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_184
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_190
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_230
timestamp 1698431365
transform 1 0 27104 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_234
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_250
timestamp 1698431365
transform 1 0 29344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_252
timestamp 1698431365
transform 1 0 29568 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_257
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_259
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_268
timestamp 1698431365
transform 1 0 31360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_272
timestamp 1698431365
transform 1 0 31808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_297
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_308
timestamp 1698431365
transform 1 0 35840 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_312
timestamp 1698431365
transform 1 0 36288 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_315
timestamp 1698431365
transform 1 0 36624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_319
timestamp 1698431365
transform 1 0 37072 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_335
timestamp 1698431365
transform 1 0 38864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_343
timestamp 1698431365
transform 1 0 39760 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_366
timestamp 1698431365
transform 1 0 42336 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_406
timestamp 1698431365
transform 1 0 46816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_410
timestamp 1698431365
transform 1 0 47264 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_434
timestamp 1698431365
transform 1 0 49952 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_450
timestamp 1698431365
transform 1 0 51744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_458
timestamp 1698431365
transform 1 0 52640 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_12
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_16
timestamp 1698431365
transform 1 0 3136 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_20
timestamp 1698431365
transform 1 0 3584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_41
timestamp 1698431365
transform 1 0 5936 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_48
timestamp 1698431365
transform 1 0 6720 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_102
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_111
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_120
timestamp 1698431365
transform 1 0 14784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_122
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_129
timestamp 1698431365
transform 1 0 15792 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_138
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_142
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_158
timestamp 1698431365
transform 1 0 19040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_162
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_196
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_202
timestamp 1698431365
transform 1 0 23968 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_206
timestamp 1698431365
transform 1 0 24416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_215
timestamp 1698431365
transform 1 0 25424 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_257
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_276
timestamp 1698431365
transform 1 0 32256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_278
timestamp 1698431365
transform 1 0 32480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_299
timestamp 1698431365
transform 1 0 34832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698431365
transform 1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_319
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_328
timestamp 1698431365
transform 1 0 38080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_330
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_349
timestamp 1698431365
transform 1 0 40432 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_365
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_395
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_411
timestamp 1698431365
transform 1 0 47376 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_427
timestamp 1698431365
transform 1 0 49168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_435
timestamp 1698431365
transform 1 0 50064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_437
timestamp 1698431365
transform 1 0 50288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_450
timestamp 1698431365
transform 1 0 51744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_461
timestamp 1698431365
transform 1 0 52976 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_477
timestamp 1698431365
transform 1 0 54768 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_481
timestamp 1698431365
transform 1 0 55216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_14
timestamp 1698431365
transform 1 0 2912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_26
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_125
timestamp 1698431365
transform 1 0 15344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698431365
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_158
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_230
timestamp 1698431365
transform 1 0 27104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_234
timestamp 1698431365
transform 1 0 27552 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_238
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_244
timestamp 1698431365
transform 1 0 28672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_248
timestamp 1698431365
transform 1 0 29120 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_266
timestamp 1698431365
transform 1 0 31136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_306
timestamp 1698431365
transform 1 0 35616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_320
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_328
timestamp 1698431365
transform 1 0 38080 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_362
timestamp 1698431365
transform 1 0 41888 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_376
timestamp 1698431365
transform 1 0 43456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_380
timestamp 1698431365
transform 1 0 43904 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_410
timestamp 1698431365
transform 1 0 47264 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_434
timestamp 1698431365
transform 1 0 49952 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_481
timestamp 1698431365
transform 1 0 55216 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_489
timestamp 1698431365
transform 1 0 56112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_61
timestamp 1698431365
transform 1 0 8176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_65
timestamp 1698431365
transform 1 0 8624 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_78
timestamp 1698431365
transform 1 0 10080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_82
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_90
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_119
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_121
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_200
timestamp 1698431365
transform 1 0 23744 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_218
timestamp 1698431365
transform 1 0 25760 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_222
timestamp 1698431365
transform 1 0 26208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_224
timestamp 1698431365
transform 1 0 26432 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_227
timestamp 1698431365
transform 1 0 26768 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_265
timestamp 1698431365
transform 1 0 31024 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_281
timestamp 1698431365
transform 1 0 32816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_295
timestamp 1698431365
transform 1 0 34384 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_361
timestamp 1698431365
transform 1 0 41776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_369
timestamp 1698431365
transform 1 0 42672 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_379
timestamp 1698431365
transform 1 0 43792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_413
timestamp 1698431365
transform 1 0 47600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_421
timestamp 1698431365
transform 1 0 48496 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_428
timestamp 1698431365
transform 1 0 49280 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_437
timestamp 1698431365
transform 1 0 50288 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_445
timestamp 1698431365
transform 1 0 51184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_452
timestamp 1698431365
transform 1 0 51968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_454
timestamp 1698431365
transform 1 0 52192 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_465
timestamp 1698431365
transform 1 0 53424 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_481
timestamp 1698431365
transform 1 0 55216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_8
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_28
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_110
timestamp 1698431365
transform 1 0 13664 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_126
timestamp 1698431365
transform 1 0 15456 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_134
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_164
timestamp 1698431365
transform 1 0 19712 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_180
timestamp 1698431365
transform 1 0 21504 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_188
timestamp 1698431365
transform 1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_190
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_197
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_203
timestamp 1698431365
transform 1 0 24080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_223
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_245
timestamp 1698431365
transform 1 0 28784 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_249
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_269
timestamp 1698431365
transform 1 0 31472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_273
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698431365
transform 1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_322
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_340
timestamp 1698431365
transform 1 0 39424 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_348
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_391
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1698431365
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_426
timestamp 1698431365
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_454
timestamp 1698431365
transform 1 0 52192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_474
timestamp 1698431365
transform 1 0 54432 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_6
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_22
timestamp 1698431365
transform 1 0 3808 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_30
timestamp 1698431365
transform 1 0 4704 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_39
timestamp 1698431365
transform 1 0 5712 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_46
timestamp 1698431365
transform 1 0 6496 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_78
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_94
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_141
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_149
timestamp 1698431365
transform 1 0 18032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_156
timestamp 1698431365
transform 1 0 18816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_160
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_200
timestamp 1698431365
transform 1 0 23744 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_204
timestamp 1698431365
transform 1 0 24192 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_207
timestamp 1698431365
transform 1 0 24528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_253
timestamp 1698431365
transform 1 0 29680 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_296
timestamp 1698431365
transform 1 0 34496 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_323
timestamp 1698431365
transform 1 0 37520 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_365
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_367
timestamp 1698431365
transform 1 0 42448 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_378
timestamp 1698431365
transform 1 0 43680 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_489
timestamp 1698431365
transform 1 0 56112 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_505
timestamp 1698431365
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_106
timestamp 1698431365
transform 1 0 13216 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698431365
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698431365
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_196
timestamp 1698431365
transform 1 0 23296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_198
timestamp 1698431365
transform 1 0 23520 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_205
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_232
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_245
timestamp 1698431365
transform 1 0 28784 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_259
timestamp 1698431365
transform 1 0 30352 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_275
timestamp 1698431365
transform 1 0 32144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_284
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_291
timestamp 1698431365
transform 1 0 33936 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_299
timestamp 1698431365
transform 1 0 34832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_344
timestamp 1698431365
transform 1 0 39872 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_348
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_356
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_358
timestamp 1698431365
transform 1 0 41440 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_393
timestamp 1698431365
transform 1 0 45360 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_409
timestamp 1698431365
transform 1 0 47152 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_417
timestamp 1698431365
transform 1 0 48048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_10
timestamp 1698431365
transform 1 0 2464 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_26
timestamp 1698431365
transform 1 0 4256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_119
timestamp 1698431365
transform 1 0 14672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_139
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_161
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_165
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_181
timestamp 1698431365
transform 1 0 21616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_189
timestamp 1698431365
transform 1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_216
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_220
timestamp 1698431365
transform 1 0 25984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_222
timestamp 1698431365
transform 1 0 26208 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_229
timestamp 1698431365
transform 1 0 26992 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_286
timestamp 1698431365
transform 1 0 33376 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_294
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_301
timestamp 1698431365
transform 1 0 35056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_303
timestamp 1698431365
transform 1 0 35280 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_333
timestamp 1698431365
transform 1 0 38640 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_340
timestamp 1698431365
transform 1 0 39424 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_372
timestamp 1698431365
transform 1 0 43008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_380
timestamp 1698431365
transform 1 0 43904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_489
timestamp 1698431365
transform 1 0 56112 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_505
timestamp 1698431365
transform 1 0 57904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_28
timestamp 1698431365
transform 1 0 4480 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_78
timestamp 1698431365
transform 1 0 10080 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_94
timestamp 1698431365
transform 1 0 11872 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_96
timestamp 1698431365
transform 1 0 12096 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_109
timestamp 1698431365
transform 1 0 13552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_113
timestamp 1698431365
transform 1 0 14000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_115
timestamp 1698431365
transform 1 0 14224 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_167
timestamp 1698431365
transform 1 0 20048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_171
timestamp 1698431365
transform 1 0 20496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_189
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_195
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_258
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_274
timestamp 1698431365
transform 1 0 32032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_316
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_324
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_328
timestamp 1698431365
transform 1 0 38080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_337
timestamp 1698431365
transform 1 0 39088 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_356
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_358
timestamp 1698431365
transform 1 0 41440 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_393
timestamp 1698431365
transform 1 0 45360 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_409
timestamp 1698431365
transform 1 0 47152 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_417
timestamp 1698431365
transform 1 0 48048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_500
timestamp 1698431365
transform 1 0 57344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_73
timestamp 1698431365
transform 1 0 9520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_75
timestamp 1698431365
transform 1 0 9744 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_111
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_121
timestamp 1698431365
transform 1 0 14896 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_153
timestamp 1698431365
transform 1 0 18480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_155
timestamp 1698431365
transform 1 0 18704 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_158
timestamp 1698431365
transform 1 0 19040 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_197
timestamp 1698431365
transform 1 0 23408 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_201
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_219
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_223
timestamp 1698431365
transform 1 0 26320 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_226
timestamp 1698431365
transform 1 0 26656 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_242
timestamp 1698431365
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_249
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_252
timestamp 1698431365
transform 1 0 29568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_284
timestamp 1698431365
transform 1 0 33152 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_300
timestamp 1698431365
transform 1 0 34944 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_308
timestamp 1698431365
transform 1 0 35840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_347
timestamp 1698431365
transform 1 0 40208 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_379
timestamp 1698431365
transform 1 0 43792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_489
timestamp 1698431365
transform 1 0 56112 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_505
timestamp 1698431365
transform 1 0 57904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_38
timestamp 1698431365
transform 1 0 5600 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_54
timestamp 1698431365
transform 1 0 7392 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_62
timestamp 1698431365
transform 1 0 8288 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_90
timestamp 1698431365
transform 1 0 11424 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_102
timestamp 1698431365
transform 1 0 12768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_104
timestamp 1698431365
transform 1 0 12992 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_131
timestamp 1698431365
transform 1 0 16016 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_168
timestamp 1698431365
transform 1 0 20160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_172
timestamp 1698431365
transform 1 0 20608 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_189
timestamp 1698431365
transform 1 0 22512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_199
timestamp 1698431365
transform 1 0 23632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_216
timestamp 1698431365
transform 1 0 25536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_236
timestamp 1698431365
transform 1 0 27776 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_239
timestamp 1698431365
transform 1 0 28112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_243
timestamp 1698431365
transform 1 0 28560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_256
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_261
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_275
timestamp 1698431365
transform 1 0 32144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_316
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_345
timestamp 1698431365
transform 1 0 39984 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_394
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_410
timestamp 1698431365
transform 1 0 47264 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_111
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_144
timestamp 1698431365
transform 1 0 17472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_164
timestamp 1698431365
transform 1 0 19712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_166
timestamp 1698431365
transform 1 0 19936 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_228
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_267
timestamp 1698431365
transform 1 0 31248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_303
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_307
timestamp 1698431365
transform 1 0 35728 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_335
timestamp 1698431365
transform 1 0 38864 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_343
timestamp 1698431365
transform 1 0 39760 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_350
timestamp 1698431365
transform 1 0 40544 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_358
timestamp 1698431365
transform 1 0 41440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_360
timestamp 1698431365
transform 1 0 41664 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_367
timestamp 1698431365
transform 1 0 42448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_374
timestamp 1698431365
transform 1 0 43232 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_393
timestamp 1698431365
transform 1 0 45360 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_425
timestamp 1698431365
transform 1 0 48944 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_441
timestamp 1698431365
transform 1 0 50736 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_449
timestamp 1698431365
transform 1 0 51632 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698431365
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_489
timestamp 1698431365
transform 1 0 56112 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_28
timestamp 1698431365
transform 1 0 4480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_32
timestamp 1698431365
transform 1 0 4928 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_48
timestamp 1698431365
transform 1 0 6720 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_56
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_60
timestamp 1698431365
transform 1 0 8064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_116
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_130
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_144
timestamp 1698431365
transform 1 0 17472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_197
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_288
timestamp 1698431365
transform 1 0 33600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_292
timestamp 1698431365
transform 1 0 34048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_294
timestamp 1698431365
transform 1 0 34272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_329
timestamp 1698431365
transform 1 0 38192 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_345
timestamp 1698431365
transform 1 0 39984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_368
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_372
timestamp 1698431365
transform 1 0 43008 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_388
timestamp 1698431365
transform 1 0 44800 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_500
timestamp 1698431365
transform 1 0 57344 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_504
timestamp 1698431365
transform 1 0 57792 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_61
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_73
timestamp 1698431365
transform 1 0 9520 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_127
timestamp 1698431365
transform 1 0 15568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_129
timestamp 1698431365
transform 1 0 15792 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_164
timestamp 1698431365
transform 1 0 19712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_168
timestamp 1698431365
transform 1 0 20160 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_207
timestamp 1698431365
transform 1 0 24528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_213
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_234
timestamp 1698431365
transform 1 0 27552 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_269
timestamp 1698431365
transform 1 0 31472 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_273
timestamp 1698431365
transform 1 0 31920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_275
timestamp 1698431365
transform 1 0 32144 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_280
timestamp 1698431365
transform 1 0 32704 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_310
timestamp 1698431365
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_341
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_343
timestamp 1698431365
transform 1 0 39760 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_359
timestamp 1698431365
transform 1 0 41552 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_375
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_473
timestamp 1698431365
transform 1 0 54320 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_481
timestamp 1698431365
transform 1 0 55216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_50
timestamp 1698431365
transform 1 0 6944 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_54
timestamp 1698431365
transform 1 0 7392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_82
timestamp 1698431365
transform 1 0 10528 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_200
timestamp 1698431365
transform 1 0 23744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_269
timestamp 1698431365
transform 1 0 31472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_273
timestamp 1698431365
transform 1 0 31920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_318
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_334
timestamp 1698431365
transform 1 0 38752 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_340
timestamp 1698431365
transform 1 0 39424 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_347
timestamp 1698431365
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_374
timestamp 1698431365
transform 1 0 43232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_387
timestamp 1698431365
transform 1 0 44688 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_395
timestamp 1698431365
transform 1 0 45584 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_399
timestamp 1698431365
transform 1 0 46032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_407
timestamp 1698431365
transform 1 0 46928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_415
timestamp 1698431365
transform 1 0 47824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_148
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_222
timestamp 1698431365
transform 1 0 26208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_233
timestamp 1698431365
transform 1 0 27440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_235
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_413
timestamp 1698431365
transform 1 0 47600 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_445
timestamp 1698431365
transform 1 0 51184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_453
timestamp 1698431365
transform 1 0 52080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_473
timestamp 1698431365
transform 1 0 54320 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_481
timestamp 1698431365
transform 1 0 55216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_34
timestamp 1698431365
transform 1 0 5152 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_50
timestamp 1698431365
transform 1 0 6944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_168
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_172
timestamp 1698431365
transform 1 0 20608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_236
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_240
timestamp 1698431365
transform 1 0 28224 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_256
timestamp 1698431365
transform 1 0 30016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_260
timestamp 1698431365
transform 1 0 30464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_273
timestamp 1698431365
transform 1 0 31920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698431365
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_288
timestamp 1698431365
transform 1 0 33600 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_307
timestamp 1698431365
transform 1 0 35728 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_315
timestamp 1698431365
transform 1 0 36624 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_334
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_336
timestamp 1698431365
transform 1 0 38976 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_348
timestamp 1698431365
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_365
timestamp 1698431365
transform 1 0 42224 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_373
timestamp 1698431365
transform 1 0 43120 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_385
timestamp 1698431365
transform 1 0 44464 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_401
timestamp 1698431365
transform 1 0 46256 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_403
timestamp 1698431365
transform 1 0 46480 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_412
timestamp 1698431365
transform 1 0 47488 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_22
timestamp 1698431365
transform 1 0 3808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_61
timestamp 1698431365
transform 1 0 8176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_65
timestamp 1698431365
transform 1 0 8624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_67
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_76
timestamp 1698431365
transform 1 0 9856 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_109
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_152
timestamp 1698431365
transform 1 0 18368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_154
timestamp 1698431365
transform 1 0 18592 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_165
timestamp 1698431365
transform 1 0 19824 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_179
timestamp 1698431365
transform 1 0 21392 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_188
timestamp 1698431365
transform 1 0 22400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_190
timestamp 1698431365
transform 1 0 22624 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_225
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_229
timestamp 1698431365
transform 1 0 26992 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_260
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_264
timestamp 1698431365
transform 1 0 30912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_268
timestamp 1698431365
transform 1 0 31360 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_307
timestamp 1698431365
transform 1 0 35728 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_328
timestamp 1698431365
transform 1 0 38080 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_360
timestamp 1698431365
transform 1 0 41664 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_364
timestamp 1698431365
transform 1 0 42112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_371
timestamp 1698431365
transform 1 0 42896 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_379
timestamp 1698431365
transform 1 0 43792 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_432
timestamp 1698431365
transform 1 0 49728 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_448
timestamp 1698431365
transform 1 0 51520 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_452
timestamp 1698431365
transform 1 0 51968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1698431365
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_473
timestamp 1698431365
transform 1 0 54320 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_481
timestamp 1698431365
transform 1 0 55216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_34
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_50
timestamp 1698431365
transform 1 0 6944 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_58
timestamp 1698431365
transform 1 0 7840 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_62
timestamp 1698431365
transform 1 0 8288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_78
timestamp 1698431365
transform 1 0 10080 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_87
timestamp 1698431365
transform 1 0 11088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_115
timestamp 1698431365
transform 1 0 14224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_148
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_164
timestamp 1698431365
transform 1 0 19712 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_183
timestamp 1698431365
transform 1 0 21840 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_272
timestamp 1698431365
transform 1 0 31808 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_289
timestamp 1698431365
transform 1 0 33712 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_299
timestamp 1698431365
transform 1 0 34832 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_331
timestamp 1698431365
transform 1 0 38416 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_339
timestamp 1698431365
transform 1 0 39312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_341
timestamp 1698431365
transform 1 0 39536 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_344
timestamp 1698431365
transform 1 0 39872 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_354
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_357
timestamp 1698431365
transform 1 0 41328 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_380
timestamp 1698431365
transform 1 0 43904 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_396
timestamp 1698431365
transform 1 0 45696 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_500
timestamp 1698431365
transform 1 0 57344 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_504
timestamp 1698431365
transform 1 0 57792 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_53
timestamp 1698431365
transform 1 0 7280 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_61
timestamp 1698431365
transform 1 0 8176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_79
timestamp 1698431365
transform 1 0 10192 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_152
timestamp 1698431365
transform 1 0 18368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_164
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_182
timestamp 1698431365
transform 1 0 21728 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_186
timestamp 1698431365
transform 1 0 22176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_188
timestamp 1698431365
transform 1 0 22400 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_261
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_300
timestamp 1698431365
transform 1 0 34944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_302
timestamp 1698431365
transform 1 0 35168 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_371
timestamp 1698431365
transform 1 0 42896 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_389
timestamp 1698431365
transform 1 0 44912 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_398
timestamp 1698431365
transform 1 0 45920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_400
timestamp 1698431365
transform 1 0 46144 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_409
timestamp 1698431365
transform 1 0 47152 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_441
timestamp 1698431365
transform 1 0 50736 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_449
timestamp 1698431365
transform 1 0 51632 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_453
timestamp 1698431365
transform 1 0 52080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_489
timestamp 1698431365
transform 1 0 56112 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_130
timestamp 1698431365
transform 1 0 15904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_132
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_163
timestamp 1698431365
transform 1 0 19600 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_342
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_383
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_415
timestamp 1698431365
transform 1 0 47824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_440
timestamp 1698431365
transform 1 0 50624 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_472
timestamp 1698431365
transform 1 0 54208 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_488
timestamp 1698431365
transform 1 0 56000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_6
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_22
timestamp 1698431365
transform 1 0 3808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_53
timestamp 1698431365
transform 1 0 7280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_61
timestamp 1698431365
transform 1 0 8176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_63
timestamp 1698431365
transform 1 0 8400 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_86
timestamp 1698431365
transform 1 0 10976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_90
timestamp 1698431365
transform 1 0 11424 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_103
timestamp 1698431365
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_126
timestamp 1698431365
transform 1 0 15456 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_130
timestamp 1698431365
transform 1 0 15904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_140
timestamp 1698431365
transform 1 0 17024 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_148
timestamp 1698431365
transform 1 0 17920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_150
timestamp 1698431365
transform 1 0 18144 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_167
timestamp 1698431365
transform 1 0 20048 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_179
timestamp 1698431365
transform 1 0 21392 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_182
timestamp 1698431365
transform 1 0 21728 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_226
timestamp 1698431365
transform 1 0 26656 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_235
timestamp 1698431365
transform 1 0 27664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_299
timestamp 1698431365
transform 1 0 34832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_303
timestamp 1698431365
transform 1 0 35280 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_343
timestamp 1698431365
transform 1 0 39760 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_375
timestamp 1698431365
transform 1 0 43344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_383
timestamp 1698431365
transform 1 0 44240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_395
timestamp 1698431365
transform 1 0 45584 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_419
timestamp 1698431365
transform 1 0 48272 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_435
timestamp 1698431365
transform 1 0 50064 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_473
timestamp 1698431365
transform 1 0 54320 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_481
timestamp 1698431365
transform 1 0 55216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_80
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_88
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_97
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_101
timestamp 1698431365
transform 1 0 12656 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_117
timestamp 1698431365
transform 1 0 14448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_121
timestamp 1698431365
transform 1 0 14896 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_146
timestamp 1698431365
transform 1 0 17696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_159
timestamp 1698431365
transform 1 0 19152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_163
timestamp 1698431365
transform 1 0 19600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_165
timestamp 1698431365
transform 1 0 19824 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_168
timestamp 1698431365
transform 1 0 20160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_176
timestamp 1698431365
transform 1 0 21056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_188
timestamp 1698431365
transform 1 0 22400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_313
timestamp 1698431365
transform 1 0 36400 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_329
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_359
timestamp 1698431365
transform 1 0 41552 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_375
timestamp 1698431365
transform 1 0 43344 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_389
timestamp 1698431365
transform 1 0 44912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_391
timestamp 1698431365
transform 1 0 45136 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_402
timestamp 1698431365
transform 1 0 46368 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_411
timestamp 1698431365
transform 1 0 47376 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_430
timestamp 1698431365
transform 1 0 49504 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_452
timestamp 1698431365
transform 1 0 51968 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_484
timestamp 1698431365
transform 1 0 55552 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_488
timestamp 1698431365
transform 1 0 56000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_73
timestamp 1698431365
transform 1 0 9520 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_75
timestamp 1698431365
transform 1 0 9744 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_84
timestamp 1698431365
transform 1 0 10752 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_90
timestamp 1698431365
transform 1 0 11424 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_98
timestamp 1698431365
transform 1 0 12320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698431365
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_134
timestamp 1698431365
transform 1 0 16352 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_138
timestamp 1698431365
transform 1 0 16800 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_159
timestamp 1698431365
transform 1 0 19152 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_161
timestamp 1698431365
transform 1 0 19376 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_191
timestamp 1698431365
transform 1 0 22736 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_195
timestamp 1698431365
transform 1 0 23184 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_210
timestamp 1698431365
transform 1 0 24864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_220
timestamp 1698431365
transform 1 0 25984 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_224
timestamp 1698431365
transform 1 0 26432 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_235
timestamp 1698431365
transform 1 0 27664 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_255
timestamp 1698431365
transform 1 0 29904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_257
timestamp 1698431365
transform 1 0 30128 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_273
timestamp 1698431365
transform 1 0 31920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_277
timestamp 1698431365
transform 1 0 32368 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_281
timestamp 1698431365
transform 1 0 32816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_285
timestamp 1698431365
transform 1 0 33264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_287
timestamp 1698431365
transform 1 0 33488 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_321
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_324
timestamp 1698431365
transform 1 0 37632 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_379
timestamp 1698431365
transform 1 0 43792 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_407
timestamp 1698431365
transform 1 0 46928 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_423
timestamp 1698431365
transform 1 0 48720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_445
timestamp 1698431365
transform 1 0 51184 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_453
timestamp 1698431365
transform 1 0 52080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_473
timestamp 1698431365
transform 1 0 54320 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_481
timestamp 1698431365
transform 1 0 55216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_76
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_101
timestamp 1698431365
transform 1 0 12656 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_105
timestamp 1698431365
transform 1 0 13104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_107
timestamp 1698431365
transform 1 0 13328 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_113
timestamp 1698431365
transform 1 0 14000 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_119
timestamp 1698431365
transform 1 0 14672 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_127
timestamp 1698431365
transform 1 0 15568 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_130
timestamp 1698431365
transform 1 0 15904 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_148
timestamp 1698431365
transform 1 0 17920 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_236
timestamp 1698431365
transform 1 0 27776 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_240
timestamp 1698431365
transform 1 0 28224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_250
timestamp 1698431365
transform 1 0 29344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_270
timestamp 1698431365
transform 1 0 31584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_274
timestamp 1698431365
transform 1 0 32032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_336
timestamp 1698431365
transform 1 0 38976 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_340
timestamp 1698431365
transform 1 0 39424 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_375
timestamp 1698431365
transform 1 0 43344 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_383
timestamp 1698431365
transform 1 0 44240 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_387
timestamp 1698431365
transform 1 0 44688 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_394
timestamp 1698431365
transform 1 0 45472 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_402
timestamp 1698431365
transform 1 0 46368 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_406
timestamp 1698431365
transform 1 0 46816 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_415
timestamp 1698431365
transform 1 0 47824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_419
timestamp 1698431365
transform 1 0 48272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_426
timestamp 1698431365
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_428
timestamp 1698431365
transform 1 0 49280 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_465
timestamp 1698431365
transform 1 0 53424 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_481
timestamp 1698431365
transform 1 0 55216 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_69
timestamp 1698431365
transform 1 0 9072 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_73
timestamp 1698431365
transform 1 0 9520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_75
timestamp 1698431365
transform 1 0 9744 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_122
timestamp 1698431365
transform 1 0 15008 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_195
timestamp 1698431365
transform 1 0 23184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_197
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_251
timestamp 1698431365
transform 1 0 29456 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_276
timestamp 1698431365
transform 1 0 32256 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_292
timestamp 1698431365
transform 1 0 34048 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_305
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_313
timestamp 1698431365
transform 1 0 36400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_323
timestamp 1698431365
transform 1 0 37520 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_327
timestamp 1698431365
transform 1 0 37968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_329
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_340
timestamp 1698431365
transform 1 0 39424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_344
timestamp 1698431365
transform 1 0 39872 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_360
timestamp 1698431365
transform 1 0 41664 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_364
timestamp 1698431365
transform 1 0 42112 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_378
timestamp 1698431365
transform 1 0 43680 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_382
timestamp 1698431365
transform 1 0 44128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_421
timestamp 1698431365
transform 1 0 48496 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_437
timestamp 1698431365
transform 1 0 50288 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_447
timestamp 1698431365
transform 1 0 51408 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_463
timestamp 1698431365
transform 1 0 53200 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_479
timestamp 1698431365
transform 1 0 54992 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_135
timestamp 1698431365
transform 1 0 16464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1698431365
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_150
timestamp 1698431365
transform 1 0 18144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_154
timestamp 1698431365
transform 1 0 18592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_158
timestamp 1698431365
transform 1 0 19040 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_162
timestamp 1698431365
transform 1 0 19488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_169
timestamp 1698431365
transform 1 0 20272 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_202
timestamp 1698431365
transform 1 0 23968 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_222
timestamp 1698431365
transform 1 0 26208 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_230
timestamp 1698431365
transform 1 0 27104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_232
timestamp 1698431365
transform 1 0 27328 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_258
timestamp 1698431365
transform 1 0 30240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_274
timestamp 1698431365
transform 1 0 32032 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_290
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_300
timestamp 1698431365
transform 1 0 34944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_304
timestamp 1698431365
transform 1 0 35392 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_320
timestamp 1698431365
transform 1 0 37184 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_324
timestamp 1698431365
transform 1 0 37632 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_348
timestamp 1698431365
transform 1 0 40320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_372
timestamp 1698431365
transform 1 0 43008 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_380
timestamp 1698431365
transform 1 0 43904 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_390
timestamp 1698431365
transform 1 0 45024 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_398
timestamp 1698431365
transform 1 0 45920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_405
timestamp 1698431365
transform 1 0 46704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_413
timestamp 1698431365
transform 1 0 47600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_417
timestamp 1698431365
transform 1 0 48048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_426
timestamp 1698431365
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_428
timestamp 1698431365
transform 1 0 49280 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_437
timestamp 1698431365
transform 1 0 50288 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_469
timestamp 1698431365
transform 1 0 53872 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_485
timestamp 1698431365
transform 1 0 55664 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698431365
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_69
timestamp 1698431365
transform 1 0 9072 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_85
timestamp 1698431365
transform 1 0 10864 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_134
timestamp 1698431365
transform 1 0 16352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_140
timestamp 1698431365
transform 1 0 17024 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_156
timestamp 1698431365
transform 1 0 18816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_160
timestamp 1698431365
transform 1 0 19264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_242
timestamp 1698431365
transform 1 0 28448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_251
timestamp 1698431365
transform 1 0 29456 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_327
timestamp 1698431365
transform 1 0 37968 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_343
timestamp 1698431365
transform 1 0 39760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_347
timestamp 1698431365
transform 1 0 40208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_351
timestamp 1698431365
transform 1 0 40656 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_367
timestamp 1698431365
transform 1 0 42448 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_375
timestamp 1698431365
transform 1 0 43344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_391
timestamp 1698431365
transform 1 0 45136 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_397
timestamp 1698431365
transform 1 0 45808 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_401
timestamp 1698431365
transform 1 0 46256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_411
timestamp 1698431365
transform 1 0 47376 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_427
timestamp 1698431365
transform 1 0 49168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_439
timestamp 1698431365
transform 1 0 50512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_443
timestamp 1698431365
transform 1 0 50960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698431365
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_464
timestamp 1698431365
transform 1 0 53312 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_496
timestamp 1698431365
transform 1 0 56896 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_504
timestamp 1698431365
transform 1 0 57792 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_508
timestamp 1698431365
transform 1 0 58240 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_80
timestamp 1698431365
transform 1 0 10304 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_84
timestamp 1698431365
transform 1 0 10752 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_86
timestamp 1698431365
transform 1 0 10976 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_95
timestamp 1698431365
transform 1 0 11984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_97
timestamp 1698431365
transform 1 0 12208 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_106
timestamp 1698431365
transform 1 0 13216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_108
timestamp 1698431365
transform 1 0 13440 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_124
timestamp 1698431365
transform 1 0 15232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_128
timestamp 1698431365
transform 1 0 15680 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_152
timestamp 1698431365
transform 1 0 18368 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_197
timestamp 1698431365
transform 1 0 23408 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698431365
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_221
timestamp 1698431365
transform 1 0 26096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_237
timestamp 1698431365
transform 1 0 27888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_241
timestamp 1698431365
transform 1 0 28336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_245
timestamp 1698431365
transform 1 0 28784 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_249
timestamp 1698431365
transform 1 0 29232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_257
timestamp 1698431365
transform 1 0 30128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_259
timestamp 1698431365
transform 1 0 30352 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_270
timestamp 1698431365
transform 1 0 31584 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_278
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_298
timestamp 1698431365
transform 1 0 34720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_306
timestamp 1698431365
transform 1 0 35616 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_338
timestamp 1698431365
transform 1 0 39200 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_359
timestamp 1698431365
transform 1 0 41552 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_394
timestamp 1698431365
transform 1 0 45472 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_396
timestamp 1698431365
transform 1 0 45696 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_438
timestamp 1698431365
transform 1 0 50400 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_472
timestamp 1698431365
transform 1 0 54208 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_488
timestamp 1698431365
transform 1 0 56000 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_69
timestamp 1698431365
transform 1 0 9072 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_85
timestamp 1698431365
transform 1 0 10864 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_93
timestamp 1698431365
transform 1 0 11760 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_97
timestamp 1698431365
transform 1 0 12208 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_100
timestamp 1698431365
transform 1 0 12544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_102
timestamp 1698431365
transform 1 0 12768 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_115
timestamp 1698431365
transform 1 0 14224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_121
timestamp 1698431365
transform 1 0 14896 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_125
timestamp 1698431365
transform 1 0 15344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_166
timestamp 1698431365
transform 1 0 19936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_168
timestamp 1698431365
transform 1 0 20160 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_174
timestamp 1698431365
transform 1 0 20832 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_179
timestamp 1698431365
transform 1 0 21392 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_182
timestamp 1698431365
transform 1 0 21728 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_186
timestamp 1698431365
transform 1 0 22176 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_211
timestamp 1698431365
transform 1 0 24976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_215
timestamp 1698431365
transform 1 0 25424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_219
timestamp 1698431365
transform 1 0 25872 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_223
timestamp 1698431365
transform 1 0 26320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_225
timestamp 1698431365
transform 1 0 26544 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_264
timestamp 1698431365
transform 1 0 30912 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_278
timestamp 1698431365
transform 1 0 32480 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_330
timestamp 1698431365
transform 1 0 38304 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_348
timestamp 1698431365
transform 1 0 40320 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_380
timestamp 1698431365
transform 1 0 43904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_384
timestamp 1698431365
transform 1 0 44352 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_391
timestamp 1698431365
transform 1 0 45136 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_397
timestamp 1698431365
transform 1 0 45808 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_401
timestamp 1698431365
transform 1 0 46256 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_409
timestamp 1698431365
transform 1 0 47152 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_425
timestamp 1698431365
transform 1 0 48944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_448
timestamp 1698431365
transform 1 0 51520 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_452
timestamp 1698431365
transform 1 0 51968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_473
timestamp 1698431365
transform 1 0 54320 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_481
timestamp 1698431365
transform 1 0 55216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_80
timestamp 1698431365
transform 1 0 10304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_84
timestamp 1698431365
transform 1 0 10752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_86
timestamp 1698431365
transform 1 0 10976 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_95
timestamp 1698431365
transform 1 0 11984 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_103
timestamp 1698431365
transform 1 0 12880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_131
timestamp 1698431365
transform 1 0 16016 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_135
timestamp 1698431365
transform 1 0 16464 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1698431365
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_150
timestamp 1698431365
transform 1 0 18144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_154
timestamp 1698431365
transform 1 0 18592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_158
timestamp 1698431365
transform 1 0 19040 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_193
timestamp 1698431365
transform 1 0 22960 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_200
timestamp 1698431365
transform 1 0 23744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_204
timestamp 1698431365
transform 1 0 24192 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_278
timestamp 1698431365
transform 1 0 32480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_296
timestamp 1698431365
transform 1 0 34496 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_309
timestamp 1698431365
transform 1 0 35952 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_325
timestamp 1698431365
transform 1 0 37744 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_356
timestamp 1698431365
transform 1 0 41216 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_360
timestamp 1698431365
transform 1 0 41664 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_362
timestamp 1698431365
transform 1 0 41888 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_371
timestamp 1698431365
transform 1 0 42896 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_398
timestamp 1698431365
transform 1 0 45920 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_414
timestamp 1698431365
transform 1 0 47712 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_418
timestamp 1698431365
transform 1 0 48160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_442
timestamp 1698431365
transform 1 0 50848 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_474
timestamp 1698431365
transform 1 0 54432 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_115
timestamp 1698431365
transform 1 0 14224 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_117
timestamp 1698431365
transform 1 0 14448 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_235
timestamp 1698431365
transform 1 0 27664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_239
timestamp 1698431365
transform 1 0 28112 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_251
timestamp 1698431365
transform 1 0 29456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_271
timestamp 1698431365
transform 1 0 31696 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_279
timestamp 1698431365
transform 1 0 32592 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_321
timestamp 1698431365
transform 1 0 37296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_323
timestamp 1698431365
transform 1 0 37520 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_326
timestamp 1698431365
transform 1 0 37856 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_334
timestamp 1698431365
transform 1 0 38752 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_350
timestamp 1698431365
transform 1 0 40544 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_358
timestamp 1698431365
transform 1 0 41440 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_360
timestamp 1698431365
transform 1 0 41664 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_395
timestamp 1698431365
transform 1 0 45584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_405
timestamp 1698431365
transform 1 0 46704 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_409
timestamp 1698431365
transform 1 0 47152 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_417
timestamp 1698431365
transform 1 0 48048 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_421
timestamp 1698431365
transform 1 0 48496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_423
timestamp 1698431365
transform 1 0 48720 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_446
timestamp 1698431365
transform 1 0 51296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_454
timestamp 1698431365
transform 1 0 52192 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_489
timestamp 1698431365
transform 1 0 56112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_80
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_84
timestamp 1698431365
transform 1 0 10752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_86
timestamp 1698431365
transform 1 0 10976 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_89
timestamp 1698431365
transform 1 0 11312 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_116
timestamp 1698431365
transform 1 0 14336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_120
timestamp 1698431365
transform 1 0 14784 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_154
timestamp 1698431365
transform 1 0 18592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_156
timestamp 1698431365
transform 1 0 18816 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_196
timestamp 1698431365
transform 1 0 23296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_231
timestamp 1698431365
transform 1 0 27216 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_235
timestamp 1698431365
transform 1 0 27664 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_245
timestamp 1698431365
transform 1 0 28784 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_268
timestamp 1698431365
transform 1 0 31360 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_290
timestamp 1698431365
transform 1 0 33824 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_297
timestamp 1698431365
transform 1 0 34608 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_301
timestamp 1698431365
transform 1 0 35056 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_330
timestamp 1698431365
transform 1 0 38304 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_338
timestamp 1698431365
transform 1 0 39200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_368
timestamp 1698431365
transform 1 0 42560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_370
timestamp 1698431365
transform 1 0 42784 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_376
timestamp 1698431365
transform 1 0 43456 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_384
timestamp 1698431365
transform 1 0 44352 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_388
timestamp 1698431365
transform 1 0 44800 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_408
timestamp 1698431365
transform 1 0 47040 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_417
timestamp 1698431365
transform 1 0 48048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1698431365
transform 1 0 48272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_430
timestamp 1698431365
transform 1 0 49504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_440
timestamp 1698431365
transform 1 0 50624 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_472
timestamp 1698431365
transform 1 0 54208 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_488
timestamp 1698431365
transform 1 0 56000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_500
timestamp 1698431365
transform 1 0 57344 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_504
timestamp 1698431365
transform 1 0 57792 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_115
timestamp 1698431365
transform 1 0 14224 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_126
timestamp 1698431365
transform 1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_130
timestamp 1698431365
transform 1 0 15904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_132
timestamp 1698431365
transform 1 0 16128 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_141
timestamp 1698431365
transform 1 0 17136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_151
timestamp 1698431365
transform 1 0 18256 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_165
timestamp 1698431365
transform 1 0 19824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_167
timestamp 1698431365
transform 1 0 20048 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_181
timestamp 1698431365
transform 1 0 21616 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_183
timestamp 1698431365
transform 1 0 21840 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_197
timestamp 1698431365
transform 1 0 23408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_205
timestamp 1698431365
transform 1 0 24304 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_209
timestamp 1698431365
transform 1 0 24752 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_217
timestamp 1698431365
transform 1 0 25648 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_221
timestamp 1698431365
transform 1 0 26096 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_223
timestamp 1698431365
transform 1 0 26320 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_226
timestamp 1698431365
transform 1 0 26656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_230
timestamp 1698431365
transform 1 0 27104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_232
timestamp 1698431365
transform 1 0 27328 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_237
timestamp 1698431365
transform 1 0 27888 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_241
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_255
timestamp 1698431365
transform 1 0 29904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_257
timestamp 1698431365
transform 1 0 30128 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_260
timestamp 1698431365
transform 1 0 30464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_273
timestamp 1698431365
transform 1 0 31920 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_286
timestamp 1698431365
transform 1 0 33376 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_302
timestamp 1698431365
transform 1 0 35168 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_310
timestamp 1698431365
transform 1 0 36064 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_341
timestamp 1698431365
transform 1 0 39536 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_345
timestamp 1698431365
transform 1 0 39984 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_361
timestamp 1698431365
transform 1 0 41776 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_369
timestamp 1698431365
transform 1 0 42672 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_377
timestamp 1698431365
transform 1 0 43568 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_379
timestamp 1698431365
transform 1 0 43792 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_399
timestamp 1698431365
transform 1 0 46032 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_426
timestamp 1698431365
transform 1 0 49056 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_434
timestamp 1698431365
transform 1 0 49952 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_436
timestamp 1698431365
transform 1 0 50176 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_450
timestamp 1698431365
transform 1 0 51744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_462
timestamp 1698431365
transform 1 0 53088 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_478
timestamp 1698431365
transform 1 0 54880 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_482
timestamp 1698431365
transform 1 0 55328 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_104
timestamp 1698431365
transform 1 0 12992 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_112
timestamp 1698431365
transform 1 0 13888 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_116
timestamp 1698431365
transform 1 0 14336 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698431365
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_146
timestamp 1698431365
transform 1 0 17696 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_150
timestamp 1698431365
transform 1 0 18144 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_153
timestamp 1698431365
transform 1 0 18480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_205
timestamp 1698431365
transform 1 0 24304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_209
timestamp 1698431365
transform 1 0 24752 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_220
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_256
timestamp 1698431365
transform 1 0 30016 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_270
timestamp 1698431365
transform 1 0 31584 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698431365
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_301
timestamp 1698431365
transform 1 0 35056 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_305
timestamp 1698431365
transform 1 0 35504 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_307
timestamp 1698431365
transform 1 0 35728 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_320
timestamp 1698431365
transform 1 0 37184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_343
timestamp 1698431365
transform 1 0 39760 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1698431365
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698431365
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_383
timestamp 1698431365
transform 1 0 44240 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_387
timestamp 1698431365
transform 1 0 44688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_402
timestamp 1698431365
transform 1 0 46368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_404
timestamp 1698431365
transform 1 0 46592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_413
timestamp 1698431365
transform 1 0 47600 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_417
timestamp 1698431365
transform 1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698431365
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_438
timestamp 1698431365
transform 1 0 50400 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_471
timestamp 1698431365
transform 1 0 54096 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_487
timestamp 1698431365
transform 1 0 55888 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1698431365
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_500
timestamp 1698431365
transform 1 0 57344 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_504
timestamp 1698431365
transform 1 0 57792 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_123
timestamp 1698431365
transform 1 0 15120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_135
timestamp 1698431365
transform 1 0 16464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_141
timestamp 1698431365
transform 1 0 17136 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_167
timestamp 1698431365
transform 1 0 20048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_169
timestamp 1698431365
transform 1 0 20272 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_223
timestamp 1698431365
transform 1 0 26320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_242
timestamp 1698431365
transform 1 0 28448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698431365
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_251
timestamp 1698431365
transform 1 0 29456 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_270
timestamp 1698431365
transform 1 0 31584 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_286
timestamp 1698431365
transform 1 0 33376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_290
timestamp 1698431365
transform 1 0 33824 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_299
timestamp 1698431365
transform 1 0 34832 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_327
timestamp 1698431365
transform 1 0 37968 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_359
timestamp 1698431365
transform 1 0 41552 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_400
timestamp 1698431365
transform 1 0 46144 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_408
timestamp 1698431365
transform 1 0 47040 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_418
timestamp 1698431365
transform 1 0 48160 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_434
timestamp 1698431365
transform 1 0 49952 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_438
timestamp 1698431365
transform 1 0 50400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_440
timestamp 1698431365
transform 1 0 50624 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_453
timestamp 1698431365
transform 1 0 52080 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698431365
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_104
timestamp 1698431365
transform 1 0 12992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_120
timestamp 1698431365
transform 1 0 14784 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_124
timestamp 1698431365
transform 1 0 15232 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_147
timestamp 1698431365
transform 1 0 17808 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_149
timestamp 1698431365
transform 1 0 18032 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_175
timestamp 1698431365
transform 1 0 20944 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_179
timestamp 1698431365
transform 1 0 21392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_181
timestamp 1698431365
transform 1 0 21616 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_194
timestamp 1698431365
transform 1 0 23072 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_198
timestamp 1698431365
transform 1 0 23520 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_208
timestamp 1698431365
transform 1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_222
timestamp 1698431365
transform 1 0 26208 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_225
timestamp 1698431365
transform 1 0 26544 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_233
timestamp 1698431365
transform 1 0 27440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_241
timestamp 1698431365
transform 1 0 28336 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_247
timestamp 1698431365
transform 1 0 29008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_251
timestamp 1698431365
transform 1 0 29456 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_259
timestamp 1698431365
transform 1 0 30352 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_261
timestamp 1698431365
transform 1 0 30576 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_284
timestamp 1698431365
transform 1 0 33152 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_306
timestamp 1698431365
transform 1 0 35616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_318
timestamp 1698431365
transform 1 0 36960 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_326
timestamp 1698431365
transform 1 0 37856 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_330
timestamp 1698431365
transform 1 0 38304 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_332
timestamp 1698431365
transform 1 0 38528 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_339
timestamp 1698431365
transform 1 0 39312 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_347
timestamp 1698431365
transform 1 0 40208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_384
timestamp 1698431365
transform 1 0 44352 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_400
timestamp 1698431365
transform 1 0 46144 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_438
timestamp 1698431365
transform 1 0 50400 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_457
timestamp 1698431365
transform 1 0 52528 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_500
timestamp 1698431365
transform 1 0 57344 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_504
timestamp 1698431365
transform 1 0 57792 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_123
timestamp 1698431365
transform 1 0 15120 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_127
timestamp 1698431365
transform 1 0 15568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_129
timestamp 1698431365
transform 1 0 15792 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_132
timestamp 1698431365
transform 1 0 16128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_149
timestamp 1698431365
transform 1 0 18032 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_157
timestamp 1698431365
transform 1 0 18928 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_167
timestamp 1698431365
transform 1 0 20048 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_205
timestamp 1698431365
transform 1 0 24304 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_222
timestamp 1698431365
transform 1 0 26208 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_226
timestamp 1698431365
transform 1 0 26656 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_231
timestamp 1698431365
transform 1 0 27216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_233
timestamp 1698431365
transform 1 0 27440 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_243
timestamp 1698431365
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_270
timestamp 1698431365
transform 1 0 31584 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_278
timestamp 1698431365
transform 1 0 32480 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_305
timestamp 1698431365
transform 1 0 35504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_330
timestamp 1698431365
transform 1 0 38304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_332
timestamp 1698431365
transform 1 0 38528 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_346
timestamp 1698431365
transform 1 0 40096 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_354
timestamp 1698431365
transform 1 0 40992 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_372
timestamp 1698431365
transform 1 0 43008 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_395
timestamp 1698431365
transform 1 0 45584 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_405
timestamp 1698431365
transform 1 0 46704 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_463
timestamp 1698431365
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_495
timestamp 1698431365
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_503
timestamp 1698431365
transform 1 0 57680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_507
timestamp 1698431365
transform 1 0 58128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_6
timestamp 1698431365
transform 1 0 2016 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_150
timestamp 1698431365
transform 1 0 18144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_202
timestamp 1698431365
transform 1 0 23968 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_214
timestamp 1698431365
transform 1 0 25312 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_234
timestamp 1698431365
transform 1 0 27552 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_286
timestamp 1698431365
transform 1 0 33376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_288
timestamp 1698431365
transform 1 0 33600 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_338
timestamp 1698431365
transform 1 0 39200 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_354
timestamp 1698431365
transform 1 0 40992 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_367
timestamp 1698431365
transform 1 0 42448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_371
timestamp 1698431365
transform 1 0 42896 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_391
timestamp 1698431365
transform 1 0 45136 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_424
timestamp 1698431365
transform 1 0 48832 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_444
timestamp 1698431365
transform 1 0 51072 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_471
timestamp 1698431365
transform 1 0 54096 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_487
timestamp 1698431365
transform 1 0 55888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_489
timestamp 1698431365
transform 1 0 56112 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_139
timestamp 1698431365
transform 1 0 16912 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_147
timestamp 1698431365
transform 1 0 17808 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_151
timestamp 1698431365
transform 1 0 18256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_153
timestamp 1698431365
transform 1 0 18480 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_156
timestamp 1698431365
transform 1 0 18816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_160
timestamp 1698431365
transform 1 0 19264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_170
timestamp 1698431365
transform 1 0 20384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_172
timestamp 1698431365
transform 1 0 20608 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_183
timestamp 1698431365
transform 1 0 21840 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_193
timestamp 1698431365
transform 1 0 22960 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_197
timestamp 1698431365
transform 1 0 23408 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_213
timestamp 1698431365
transform 1 0 25200 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_215
timestamp 1698431365
transform 1 0 25424 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_221
timestamp 1698431365
transform 1 0 26096 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_228
timestamp 1698431365
transform 1 0 26880 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_232
timestamp 1698431365
transform 1 0 27328 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_268
timestamp 1698431365
transform 1 0 31360 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_276
timestamp 1698431365
transform 1 0 32256 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_308
timestamp 1698431365
transform 1 0 35840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_312
timestamp 1698431365
transform 1 0 36288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_327
timestamp 1698431365
transform 1 0 37968 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_331
timestamp 1698431365
transform 1 0 38416 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_356
timestamp 1698431365
transform 1 0 41216 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_360
timestamp 1698431365
transform 1 0 41664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_370
timestamp 1698431365
transform 1 0 42784 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_378
timestamp 1698431365
transform 1 0 43680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_382
timestamp 1698431365
transform 1 0 44128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_384
timestamp 1698431365
transform 1 0 44352 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_397
timestamp 1698431365
transform 1 0 45808 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_401
timestamp 1698431365
transform 1 0 46256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_403
timestamp 1698431365
transform 1 0 46480 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_420
timestamp 1698431365
transform 1 0 48384 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_453
timestamp 1698431365
transform 1 0 52080 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_483
timestamp 1698431365
transform 1 0 55440 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_499
timestamp 1698431365
transform 1 0 57232 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_52
timestamp 1698431365
transform 1 0 7168 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_60
timestamp 1698431365
transform 1 0 8064 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_65
timestamp 1698431365
transform 1 0 8624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_67
timestamp 1698431365
transform 1 0 8848 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_78
timestamp 1698431365
transform 1 0 10080 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_83
timestamp 1698431365
transform 1 0 10640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_89
timestamp 1698431365
transform 1 0 11312 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_97
timestamp 1698431365
transform 1 0 12208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_101
timestamp 1698431365
transform 1 0 12656 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_108
timestamp 1698431365
transform 1 0 13440 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_113
timestamp 1698431365
transform 1 0 14000 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_129
timestamp 1698431365
transform 1 0 15792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_133
timestamp 1698431365
transform 1 0 16240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_135
timestamp 1698431365
transform 1 0 16464 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_154
timestamp 1698431365
transform 1 0 18592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_160
timestamp 1698431365
transform 1 0 19264 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_168
timestamp 1698431365
transform 1 0 20160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_210
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_216
timestamp 1698431365
transform 1 0 25536 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_220
timestamp 1698431365
transform 1 0 25984 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_230
timestamp 1698431365
transform 1 0 27104 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_244
timestamp 1698431365
transform 1 0 28672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_274
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_278
timestamp 1698431365
transform 1 0 32480 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_284
timestamp 1698431365
transform 1 0 33152 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_301
timestamp 1698431365
transform 1 0 35056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_305
timestamp 1698431365
transform 1 0 35504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_308
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_414
timestamp 1698431365
transform 1 0 47712 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698431365
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_474
timestamp 1698431365
transform 1 0 54432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_490
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_498
timestamp 1698431365
transform 1 0 57120 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_502
timestamp 1698431365
transform 1 0 57568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_504
timestamp 1698431365
transform 1 0 57792 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 58352 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_71 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_72
timestamp 1698431365
transform -1 0 2016 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_73
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_74
timestamp 1698431365
transform -1 0 2016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_75
timestamp 1698431365
transform 1 0 57456 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_76
timestamp 1698431365
transform 1 0 57456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_77
timestamp 1698431365
transform 1 0 57904 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_78
timestamp 1698431365
transform -1 0 2464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_79
timestamp 1698431365
transform -1 0 54432 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_80
timestamp 1698431365
transform 1 0 57904 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_81
timestamp 1698431365
transform -1 0 2016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_82
timestamp 1698431365
transform -1 0 5936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_83
timestamp 1698431365
transform 1 0 57904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_84
timestamp 1698431365
transform 1 0 57904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_85
timestamp 1698431365
transform -1 0 2016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_86
timestamp 1698431365
transform 1 0 57904 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_87
timestamp 1698431365
transform -1 0 10640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_88
timestamp 1698431365
transform 1 0 57904 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_89
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_90
timestamp 1698431365
transform -1 0 14000 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_91
timestamp 1698431365
transform 1 0 57904 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_92
timestamp 1698431365
transform -1 0 2016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_93
timestamp 1698431365
transform 1 0 57904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_94
timestamp 1698431365
transform -1 0 11312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_95
timestamp 1698431365
transform -1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_96
timestamp 1698431365
transform -1 0 2016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_97
timestamp 1698431365
transform 1 0 57904 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_98
timestamp 1698431365
transform -1 0 55328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  OQPSK_RCOSINE_ALL_99
timestamp 1698431365
transform -1 0 7952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_100 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 57904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_101
timestamp 1698431365
transform -1 0 56224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_102
timestamp 1698431365
transform -1 0 2016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_103
timestamp 1698431365
transform 1 0 57904 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_104
timestamp 1698431365
transform -1 0 8624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_105
timestamp 1698431365
transform 1 0 57904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_106
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_107
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  OQPSK_RCOSINE_ALL_108
timestamp 1698431365
transform -1 0 2016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 55440 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform 1 0 47824 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform 1 0 48496 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform 1 0 55440 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 55440 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform 1 0 55440 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 55440 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform 1 0 55440 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform 1 0 55440 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform 1 0 55440 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 51184 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 40320 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 55440 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 55440 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 55440 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 43792 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 51744 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 55440 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform 1 0 55440 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 55440 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1698431365
transform 1 0 55440 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1698431365
transform 1 0 55440 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1698431365
transform 1 0 53312 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1698431365
transform -1 0 4480 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output33
timestamp 1698431365
transform -1 0 4480 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output34
timestamp 1698431365
transform -1 0 4480 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output35
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36
timestamp 1698431365
transform -1 0 4480 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1698431365
transform -1 0 31808 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1698431365
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698431365
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698431365
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1698431365
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698431365
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
<< labels >>
flabel metal3 s 59200 30240 60000 30352 0 FreeSans 448 0 0 0 ACK
port 0 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 Bit_In
port 1 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 EN
port 2 nsew signal input
flabel metal3 s 59200 36288 60000 36400 0 FreeSans 448 0 0 0 I[0]
port 3 nsew signal tristate
flabel metal2 s 47712 59200 47824 60000 0 FreeSans 448 90 0 0 I[10]
port 4 nsew signal tristate
flabel metal2 s 49056 59200 49168 60000 0 FreeSans 448 90 0 0 I[11]
port 5 nsew signal tristate
flabel metal2 s 48384 59200 48496 60000 0 FreeSans 448 90 0 0 I[12]
port 6 nsew signal tristate
flabel metal3 s 59200 35616 60000 35728 0 FreeSans 448 0 0 0 I[1]
port 7 nsew signal tristate
flabel metal3 s 59200 37632 60000 37744 0 FreeSans 448 0 0 0 I[2]
port 8 nsew signal tristate
flabel metal3 s 59200 40320 60000 40432 0 FreeSans 448 0 0 0 I[3]
port 9 nsew signal tristate
flabel metal3 s 59200 41664 60000 41776 0 FreeSans 448 0 0 0 I[4]
port 10 nsew signal tristate
flabel metal3 s 59200 43680 60000 43792 0 FreeSans 448 0 0 0 I[5]
port 11 nsew signal tristate
flabel metal3 s 59200 47040 60000 47152 0 FreeSans 448 0 0 0 I[6]
port 12 nsew signal tristate
flabel metal3 s 59200 51072 60000 51184 0 FreeSans 448 0 0 0 I[7]
port 13 nsew signal tristate
flabel metal2 s 52416 59200 52528 60000 0 FreeSans 448 90 0 0 I[8]
port 14 nsew signal tristate
flabel metal2 s 51072 59200 51184 60000 0 FreeSans 448 90 0 0 I[9]
port 15 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 Q[0]
port 16 nsew signal tristate
flabel metal3 s 59200 26208 60000 26320 0 FreeSans 448 0 0 0 Q[10]
port 17 nsew signal tristate
flabel metal3 s 59200 27552 60000 27664 0 FreeSans 448 0 0 0 Q[11]
port 18 nsew signal tristate
flabel metal3 s 59200 24864 60000 24976 0 FreeSans 448 0 0 0 Q[12]
port 19 nsew signal tristate
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal2 s 51744 0 51856 800 0 FreeSans 448 90 0 0 Q[3]
port 22 nsew signal tristate
flabel metal3 s 59200 8736 60000 8848 0 FreeSans 448 0 0 0 Q[4]
port 23 nsew signal tristate
flabel metal3 s 59200 12096 60000 12208 0 FreeSans 448 0 0 0 Q[5]
port 24 nsew signal tristate
flabel metal3 s 59200 14784 60000 14896 0 FreeSans 448 0 0 0 Q[6]
port 25 nsew signal tristate
flabel metal3 s 59200 17472 60000 17584 0 FreeSans 448 0 0 0 Q[7]
port 26 nsew signal tristate
flabel metal3 s 59200 20832 60000 20944 0 FreeSans 448 0 0 0 Q[8]
port 27 nsew signal tristate
flabel metal3 s 59200 24192 60000 24304 0 FreeSans 448 0 0 0 Q[9]
port 28 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 REQ_SAMPLE
port 29 nsew signal input
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 RST
port 30 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 addI[0]
port 31 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 addI[1]
port 32 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 addI[2]
port 33 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 addI[3]
port 34 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 addI[4]
port 35 nsew signal tristate
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 addI[5]
port 36 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 addQ[0]
port 37 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 addQ[1]
port 38 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 addQ[2]
port 39 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 addQ[3]
port 40 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 addQ[4]
port 41 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 addQ[5]
port 42 nsew signal tristate
flabel metal3 s 59200 48384 60000 48496 0 FreeSans 448 0 0 0 io_oeb[0]
port 43 nsew signal tristate
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 io_oeb[10]
port 44 nsew signal tristate
flabel metal3 s 59200 54432 60000 54544 0 FreeSans 448 0 0 0 io_oeb[11]
port 45 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 io_oeb[12]
port 46 nsew signal tristate
flabel metal3 s 59200 55104 60000 55216 0 FreeSans 448 0 0 0 io_oeb[13]
port 47 nsew signal tristate
flabel metal3 s 59200 2688 60000 2800 0 FreeSans 448 0 0 0 io_oeb[14]
port 48 nsew signal tristate
flabel metal3 s 59200 49728 60000 49840 0 FreeSans 448 0 0 0 io_oeb[15]
port 49 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 io_oeb[16]
port 50 nsew signal tristate
flabel metal2 s 53088 59200 53200 60000 0 FreeSans 448 90 0 0 io_oeb[17]
port 51 nsew signal tristate
flabel metal3 s 59200 38304 60000 38416 0 FreeSans 448 0 0 0 io_oeb[18]
port 52 nsew signal tristate
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 io_oeb[19]
port 53 nsew signal tristate
flabel metal2 s 55104 59200 55216 60000 0 FreeSans 448 90 0 0 io_oeb[1]
port 54 nsew signal tristate
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 io_oeb[20]
port 55 nsew signal tristate
flabel metal3 s 59200 38976 60000 39088 0 FreeSans 448 0 0 0 io_oeb[21]
port 56 nsew signal tristate
flabel metal3 s 59200 32928 60000 33040 0 FreeSans 448 0 0 0 io_oeb[22]
port 57 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 io_oeb[23]
port 58 nsew signal tristate
flabel metal3 s 59200 4032 60000 4144 0 FreeSans 448 0 0 0 io_oeb[24]
port 59 nsew signal tristate
flabel metal2 s 10080 59200 10192 60000 0 FreeSans 448 90 0 0 io_oeb[25]
port 60 nsew signal tristate
flabel metal3 s 59200 33600 60000 33712 0 FreeSans 448 0 0 0 io_oeb[26]
port 61 nsew signal tristate
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_oeb[27]
port 62 nsew signal tristate
flabel metal2 s 13440 59200 13552 60000 0 FreeSans 448 90 0 0 io_oeb[28]
port 63 nsew signal tristate
flabel metal3 s 59200 49056 60000 49168 0 FreeSans 448 0 0 0 io_oeb[29]
port 64 nsew signal tristate
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 io_oeb[2]
port 65 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 io_oeb[30]
port 66 nsew signal tristate
flabel metal3 s 59200 3360 60000 3472 0 FreeSans 448 0 0 0 io_oeb[31]
port 67 nsew signal tristate
flabel metal2 s 10752 59200 10864 60000 0 FreeSans 448 90 0 0 io_oeb[32]
port 68 nsew signal tristate
flabel metal2 s 54432 59200 54544 60000 0 FreeSans 448 90 0 0 io_oeb[33]
port 69 nsew signal tristate
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 io_oeb[34]
port 70 nsew signal tristate
flabel metal3 s 59200 52416 60000 52528 0 FreeSans 448 0 0 0 io_oeb[35]
port 71 nsew signal tristate
flabel metal2 s 53760 59200 53872 60000 0 FreeSans 448 90 0 0 io_oeb[36]
port 72 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 io_oeb[37]
port 73 nsew signal tristate
flabel metal3 s 59200 55776 60000 55888 0 FreeSans 448 0 0 0 io_oeb[3]
port 74 nsew signal tristate
flabel metal2 s 8064 59200 8176 60000 0 FreeSans 448 90 0 0 io_oeb[4]
port 75 nsew signal tristate
flabel metal3 s 59200 5376 60000 5488 0 FreeSans 448 0 0 0 io_oeb[5]
port 76 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 io_oeb[6]
port 77 nsew signal tristate
flabel metal3 s 59200 4704 60000 4816 0 FreeSans 448 0 0 0 io_oeb[7]
port 78 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 io_oeb[8]
port 79 nsew signal tristate
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 io_oeb[9]
port 80 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 81 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 81 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 82 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 82 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 58184 30632 58184 30632 0 ACK
rlabel metal2 1736 26656 1736 26656 0 Bit_In
rlabel metal2 1736 27720 1736 27720 0 EN
rlabel metal2 57848 35672 57848 35672 0 I[0]
rlabel metal2 47768 57778 47768 57778 0 I[10]
rlabel metal2 49112 57778 49112 57778 0 I[11]
rlabel metal3 49056 55384 49056 55384 0 I[12]
rlabel metal2 57960 36120 57960 36120 0 I[1]
rlabel metal2 57960 37912 57960 37912 0 I[2]
rlabel metal2 57960 40824 57960 40824 0 I[3]
rlabel metal2 57960 42280 57960 42280 0 I[4]
rlabel metal2 57960 44072 57960 44072 0 I[5]
rlabel metal2 57960 47320 57960 47320 0 I[6]
rlabel metal2 57960 50960 57960 50960 0 I[7]
rlabel metal3 53088 55384 53088 55384 0 I[8]
rlabel metal3 51744 54824 51744 54824 0 I[9]
rlabel metal2 41048 2030 41048 2030 0 Q[0]
rlabel metal2 57960 25984 57960 25984 0 Q[10]
rlabel metal2 57960 27440 57960 27440 0 Q[11]
rlabel metal2 57960 24528 57960 24528 0 Q[12]
rlabel metal3 44352 3416 44352 3416 0 Q[1]
rlabel metal2 48440 1190 48440 1190 0 Q[2]
rlabel metal2 51800 2198 51800 2198 0 Q[3]
rlabel metal3 58632 8344 58632 8344 0 Q[4]
rlabel metal2 57960 12600 57960 12600 0 Q[5]
rlabel metal2 57960 14784 57960 14784 0 Q[6]
rlabel metal2 57960 17640 57960 17640 0 Q[7]
rlabel metal3 58618 20888 58618 20888 0 Q[8]
rlabel metal2 55384 24360 55384 24360 0 Q[9]
rlabel metal2 1736 25144 1736 25144 0 REQ_SAMPLE
rlabel metal2 2408 25928 2408 25928 0 RST
rlabel metal2 38248 31780 38248 31780 0 _0000_
rlabel metal2 38920 27496 38920 27496 0 _0002_
rlabel metal2 42168 33264 42168 33264 0 _0004_
rlabel metal2 31304 28728 31304 28728 0 _0005_
rlabel metal2 42616 29008 42616 29008 0 _0006_
rlabel metal2 44968 22792 44968 22792 0 _0007_
rlabel metal2 12936 28560 12936 28560 0 _0008_
rlabel metal3 15064 30184 15064 30184 0 _0009_
rlabel metal3 12152 30968 12152 30968 0 _0010_
rlabel metal2 20664 28952 20664 28952 0 _0011_
rlabel metal2 25312 28616 25312 28616 0 _0012_
rlabel metal2 26824 30688 26824 30688 0 _0013_
rlabel metal2 5600 23800 5600 23800 0 _0014_
rlabel metal3 7252 27832 7252 27832 0 _0015_
rlabel metal2 6216 25816 6216 25816 0 _0016_
rlabel metal2 9240 25928 9240 25928 0 _0017_
rlabel metal2 11816 26544 11816 26544 0 _0018_
rlabel metal3 20608 27048 20608 27048 0 _0019_
rlabel metal2 42336 30968 42336 30968 0 _0020_
rlabel metal2 42280 32928 42280 32928 0 _0021_
rlabel metal2 34328 40880 34328 40880 0 _0022_
rlabel metal3 35728 38584 35728 38584 0 _0023_
rlabel metal2 37520 37464 37520 37464 0 _0024_
rlabel metal2 39816 37296 39816 37296 0 _0025_
rlabel metal2 33600 52920 33600 52920 0 _0026_
rlabel metal3 35280 35896 35280 35896 0 _0027_
rlabel metal2 14168 36120 14168 36120 0 _0028_
rlabel metal2 13720 37072 13720 37072 0 _0029_
rlabel metal3 17696 37240 17696 37240 0 _0030_
rlabel metal3 30520 37128 30520 37128 0 _0031_
rlabel metal2 11144 36008 11144 36008 0 _0032_
rlabel metal2 31304 36232 31304 36232 0 _0033_
rlabel metal2 29848 35336 29848 35336 0 _0034_
rlabel metal2 30632 36064 30632 36064 0 _0035_
rlabel metal2 31416 36400 31416 36400 0 _0036_
rlabel metal2 35560 36120 35560 36120 0 _0037_
rlabel metal2 36904 36176 36904 36176 0 _0038_
rlabel metal2 40152 36736 40152 36736 0 _0039_
rlabel metal2 45864 36400 45864 36400 0 _0040_
rlabel metal2 45192 46144 45192 46144 0 _0041_
rlabel metal2 44408 36960 44408 36960 0 _0042_
rlabel metal2 27944 37352 27944 37352 0 _0043_
rlabel metal3 44744 36568 44744 36568 0 _0044_
rlabel metal2 47544 38780 47544 38780 0 _0045_
rlabel metal3 40264 37240 40264 37240 0 _0046_
rlabel metal3 40936 37128 40936 37128 0 _0047_
rlabel metal2 46928 39592 46928 39592 0 _0048_
rlabel metal3 40488 34104 40488 34104 0 _0049_
rlabel metal2 41272 40264 41272 40264 0 _0050_
rlabel metal2 18816 47432 18816 47432 0 _0051_
rlabel metal2 19656 44128 19656 44128 0 _0052_
rlabel metal2 16520 45976 16520 45976 0 _0053_
rlabel metal2 31080 51016 31080 51016 0 _0054_
rlabel metal2 20328 46704 20328 46704 0 _0055_
rlabel metal2 19768 41608 19768 41608 0 _0056_
rlabel metal3 8260 34664 8260 34664 0 _0057_
rlabel metal2 19096 46984 19096 46984 0 _0058_
rlabel metal2 19432 48216 19432 48216 0 _0059_
rlabel metal2 19544 46424 19544 46424 0 _0060_
rlabel metal2 28728 41888 28728 41888 0 _0061_
rlabel metal2 31752 42448 31752 42448 0 _0062_
rlabel metal2 15176 41048 15176 41048 0 _0063_
rlabel metal2 20440 38724 20440 38724 0 _0064_
rlabel metal2 29400 33040 29400 33040 0 _0065_
rlabel metal2 21672 39704 21672 39704 0 _0066_
rlabel metal3 28336 50456 28336 50456 0 _0067_
rlabel metal4 25592 49336 25592 49336 0 _0068_
rlabel metal2 27944 42056 27944 42056 0 _0069_
rlabel metal2 39592 40656 39592 40656 0 _0070_
rlabel metal3 41216 41720 41216 41720 0 _0071_
rlabel metal2 43400 39928 43400 39928 0 _0072_
rlabel metal2 35616 41048 35616 41048 0 _0073_
rlabel metal2 36568 40544 36568 40544 0 _0074_
rlabel metal2 26096 47208 26096 47208 0 _0075_
rlabel metal2 29176 34048 29176 34048 0 _0076_
rlabel metal2 26656 40264 26656 40264 0 _0077_
rlabel metal2 19208 42056 19208 42056 0 _0078_
rlabel metal3 20216 42504 20216 42504 0 _0079_
rlabel metal2 15512 43568 15512 43568 0 _0080_
rlabel metal2 8904 41496 8904 41496 0 _0081_
rlabel metal2 14952 42728 14952 42728 0 _0082_
rlabel metal2 16184 42000 16184 42000 0 _0083_
rlabel metal2 26152 42336 26152 42336 0 _0084_
rlabel metal2 26712 41776 26712 41776 0 _0085_
rlabel metal3 35112 42840 35112 42840 0 _0086_
rlabel metal2 29848 33712 29848 33712 0 _0087_
rlabel metal3 35280 37128 35280 37128 0 _0088_
rlabel metal2 23856 50120 23856 50120 0 _0089_
rlabel metal2 20104 36456 20104 36456 0 _0090_
rlabel metal3 19768 36680 19768 36680 0 _0091_
rlabel metal2 21560 36792 21560 36792 0 _0092_
rlabel metal3 19768 35560 19768 35560 0 _0093_
rlabel metal3 14868 35896 14868 35896 0 _0094_
rlabel metal3 22680 36456 22680 36456 0 _0095_
rlabel metal2 33768 37184 33768 37184 0 _0096_
rlabel metal2 34384 37240 34384 37240 0 _0097_
rlabel metal2 31192 36288 31192 36288 0 _0098_
rlabel metal2 35672 37632 35672 37632 0 _0099_
rlabel metal2 34328 37520 34328 37520 0 _0100_
rlabel metal2 37576 40096 37576 40096 0 _0101_
rlabel metal2 43512 39704 43512 39704 0 _0102_
rlabel metal3 44688 39592 44688 39592 0 _0103_
rlabel metal2 46536 38752 46536 38752 0 _0104_
rlabel metal2 47376 37464 47376 37464 0 _0105_
rlabel metal2 49056 37912 49056 37912 0 _0106_
rlabel metal3 33824 48440 33824 48440 0 _0107_
rlabel metal3 46928 38808 46928 38808 0 _0108_
rlabel metal2 46872 39088 46872 39088 0 _0109_
rlabel metal3 48496 40376 48496 40376 0 _0110_
rlabel metal2 37240 39536 37240 39536 0 _0111_
rlabel metal3 41328 39480 41328 39480 0 _0112_
rlabel metal2 46424 41216 46424 41216 0 _0113_
rlabel metal2 40040 42616 40040 42616 0 _0114_
rlabel metal3 40992 42728 40992 42728 0 _0115_
rlabel metal2 22232 44856 22232 44856 0 _0116_
rlabel metal2 23800 53872 23800 53872 0 _0117_
rlabel metal2 30968 35840 30968 35840 0 _0118_
rlabel metal2 22120 44128 22120 44128 0 _0119_
rlabel metal2 15960 45080 15960 45080 0 _0120_
rlabel metal2 20552 43792 20552 43792 0 _0121_
rlabel metal2 28616 44016 28616 44016 0 _0122_
rlabel metal3 17136 43624 17136 43624 0 _0123_
rlabel metal3 17136 44072 17136 44072 0 _0124_
rlabel metal2 20216 44240 20216 44240 0 _0125_
rlabel metal2 21784 43568 21784 43568 0 _0126_
rlabel metal2 42896 42616 42896 42616 0 _0127_
rlabel metal2 44968 43176 44968 43176 0 _0128_
rlabel metal2 13384 31556 13384 31556 0 _0129_
rlabel metal2 41496 34664 41496 34664 0 _0130_
rlabel metal2 42392 43848 42392 43848 0 _0131_
rlabel metal3 44240 43288 44240 43288 0 _0132_
rlabel metal2 45192 42336 45192 42336 0 _0133_
rlabel metal2 14168 46144 14168 46144 0 _0134_
rlabel metal2 16912 45864 16912 45864 0 _0135_
rlabel metal3 14616 45864 14616 45864 0 _0136_
rlabel metal2 16072 45864 16072 45864 0 _0137_
rlabel metal2 22512 46648 22512 46648 0 _0138_
rlabel metal2 21448 41776 21448 41776 0 _0139_
rlabel metal2 12152 31780 12152 31780 0 _0140_
rlabel metal3 16576 46760 16576 46760 0 _0141_
rlabel metal2 21784 46648 21784 46648 0 _0142_
rlabel metal2 23128 46424 23128 46424 0 _0143_
rlabel metal2 11592 45584 11592 45584 0 _0144_
rlabel metal2 23128 45304 23128 45304 0 _0145_
rlabel metal2 34328 44072 34328 44072 0 _0146_
rlabel metal2 35224 42504 35224 42504 0 _0147_
rlabel metal2 43848 42224 43848 42224 0 _0148_
rlabel metal2 20440 49056 20440 49056 0 _0149_
rlabel metal3 17136 40488 17136 40488 0 _0150_
rlabel metal3 16744 34328 16744 34328 0 _0151_
rlabel metal3 19488 39592 19488 39592 0 _0152_
rlabel metal2 20104 40572 20104 40572 0 _0153_
rlabel metal2 20720 40936 20720 40936 0 _0154_
rlabel metal2 20216 39928 20216 39928 0 _0155_
rlabel metal2 31640 37800 31640 37800 0 _0156_
rlabel metal2 21000 41720 21000 41720 0 _0157_
rlabel metal2 24864 42952 24864 42952 0 _0158_
rlabel metal2 22344 40824 22344 40824 0 _0159_
rlabel metal3 24080 38024 24080 38024 0 _0160_
rlabel metal3 25704 38024 25704 38024 0 _0161_
rlabel metal2 19544 39144 19544 39144 0 _0162_
rlabel metal2 24752 35000 24752 35000 0 _0163_
rlabel metal2 25032 35728 25032 35728 0 _0164_
rlabel metal2 31640 38080 31640 38080 0 _0165_
rlabel metal3 32984 37912 32984 37912 0 _0166_
rlabel metal3 34832 38024 34832 38024 0 _0167_
rlabel metal3 38584 37912 38584 37912 0 _0168_
rlabel metal2 43960 41216 43960 41216 0 _0169_
rlabel metal3 46648 41720 46648 41720 0 _0170_
rlabel metal2 49560 40824 49560 40824 0 _0171_
rlabel metal2 49952 40376 49952 40376 0 _0172_
rlabel metal2 28392 34720 28392 34720 0 _0173_
rlabel metal2 25928 48272 25928 48272 0 _0174_
rlabel metal2 27272 44632 27272 44632 0 _0175_
rlabel metal2 25704 46536 25704 46536 0 _0176_
rlabel metal2 27944 45752 27944 45752 0 _0177_
rlabel metal2 30128 45192 30128 45192 0 _0178_
rlabel metal2 27664 53480 27664 53480 0 _0179_
rlabel metal2 19320 49168 19320 49168 0 _0180_
rlabel metal2 25256 49728 25256 49728 0 _0181_
rlabel metal2 27048 51800 27048 51800 0 _0182_
rlabel metal2 26824 41832 26824 41832 0 _0183_
rlabel metal2 23240 51240 23240 51240 0 _0184_
rlabel metal2 29008 45192 29008 45192 0 _0185_
rlabel metal2 15064 44296 15064 44296 0 _0186_
rlabel metal4 15848 50064 15848 50064 0 _0187_
rlabel metal2 38808 44912 38808 44912 0 _0188_
rlabel metal2 39144 45136 39144 45136 0 _0189_
rlabel metal2 38416 45080 38416 45080 0 _0190_
rlabel metal3 40880 45080 40880 45080 0 _0191_
rlabel metal2 40600 51744 40600 51744 0 _0192_
rlabel metal2 47432 44632 47432 44632 0 _0193_
rlabel metal2 24136 47936 24136 47936 0 _0194_
rlabel metal2 34776 42056 34776 42056 0 _0195_
rlabel metal2 36344 43120 36344 43120 0 _0196_
rlabel metal2 25256 51072 25256 51072 0 _0197_
rlabel metal2 16184 48216 16184 48216 0 _0198_
rlabel metal2 20216 48552 20216 48552 0 _0199_
rlabel metal3 18312 45864 18312 45864 0 _0200_
rlabel metal2 18984 50232 18984 50232 0 _0201_
rlabel metal2 14168 51408 14168 51408 0 _0202_
rlabel metal2 16968 50512 16968 50512 0 _0203_
rlabel metal2 19208 52416 19208 52416 0 _0204_
rlabel metal2 30800 37800 30800 37800 0 _0205_
rlabel metal2 23464 52808 23464 52808 0 _0206_
rlabel metal2 17416 46032 17416 46032 0 _0207_
rlabel metal2 18928 50568 18928 50568 0 _0208_
rlabel metal2 19208 49616 19208 49616 0 _0209_
rlabel metal2 33768 43624 33768 43624 0 _0210_
rlabel metal3 42392 44296 42392 44296 0 _0211_
rlabel metal2 37128 50456 37128 50456 0 _0212_
rlabel metal2 34328 38360 34328 38360 0 _0213_
rlabel metal2 34440 39816 34440 39816 0 _0214_
rlabel metal2 17528 45920 17528 45920 0 _0215_
rlabel metal2 30408 36568 30408 36568 0 _0216_
rlabel metal2 17640 46592 17640 46592 0 _0217_
rlabel metal3 26852 44968 26852 44968 0 _0218_
rlabel metal3 29792 44856 29792 44856 0 _0219_
rlabel metal2 34888 44744 34888 44744 0 _0220_
rlabel metal3 36176 44296 36176 44296 0 _0221_
rlabel metal2 46200 44464 46200 44464 0 _0222_
rlabel metal2 47544 44352 47544 44352 0 _0223_
rlabel metal3 49056 43624 49056 43624 0 _0224_
rlabel metal2 45416 41440 45416 41440 0 _0225_
rlabel metal3 45304 48216 45304 48216 0 _0226_
rlabel metal2 30408 41944 30408 41944 0 _0227_
rlabel metal2 46312 42336 46312 42336 0 _0228_
rlabel metal2 49224 42448 49224 42448 0 _0229_
rlabel metal2 50792 43176 50792 43176 0 _0230_
rlabel metal2 45864 42728 45864 42728 0 _0231_
rlabel metal2 48440 41552 48440 41552 0 _0232_
rlabel metal2 50456 42560 50456 42560 0 _0233_
rlabel metal2 51296 41944 51296 41944 0 _0234_
rlabel metal2 47040 43512 47040 43512 0 _0235_
rlabel metal2 49560 44856 49560 44856 0 _0236_
rlabel metal2 30856 43904 30856 43904 0 _0237_
rlabel metal3 43288 48328 43288 48328 0 _0238_
rlabel metal2 8344 30772 8344 30772 0 _0239_
rlabel metal2 31304 51408 31304 51408 0 _0240_
rlabel metal2 25480 49336 25480 49336 0 _0241_
rlabel metal2 21336 48888 21336 48888 0 _0242_
rlabel metal2 22456 49896 22456 49896 0 _0243_
rlabel metal2 21224 54768 21224 54768 0 _0244_
rlabel metal2 13160 49840 13160 49840 0 _0245_
rlabel metal2 13608 50064 13608 50064 0 _0246_
rlabel metal2 20216 49672 20216 49672 0 _0247_
rlabel metal2 30296 49000 30296 49000 0 _0248_
rlabel metal3 21392 50456 21392 50456 0 _0249_
rlabel metal2 23296 50344 23296 50344 0 _0250_
rlabel metal2 23800 49280 23800 49280 0 _0251_
rlabel metal2 26488 48664 26488 48664 0 _0252_
rlabel metal3 41608 45752 41608 45752 0 _0253_
rlabel metal3 45360 45864 45360 45864 0 _0254_
rlabel metal2 36232 45360 36232 45360 0 _0255_
rlabel metal3 36904 47432 36904 47432 0 _0256_
rlabel metal2 30968 46396 30968 46396 0 _0257_
rlabel metal3 28672 47544 28672 47544 0 _0258_
rlabel metal2 10920 43904 10920 43904 0 _0259_
rlabel metal2 23016 47712 23016 47712 0 _0260_
rlabel metal3 23800 46928 23800 46928 0 _0261_
rlabel metal3 28728 47432 28728 47432 0 _0262_
rlabel metal2 34328 47824 34328 47824 0 _0263_
rlabel metal3 41832 47320 41832 47320 0 _0264_
rlabel metal2 46088 46480 46088 46480 0 _0265_
rlabel metal2 29232 44408 29232 44408 0 _0266_
rlabel metal2 29792 42952 29792 42952 0 _0267_
rlabel metal2 24920 42000 24920 42000 0 _0268_
rlabel metal2 31304 44016 31304 44016 0 _0269_
rlabel metal2 8680 39592 8680 39592 0 _0270_
rlabel metal2 30240 49784 30240 49784 0 _0271_
rlabel metal2 29848 47040 29848 47040 0 _0272_
rlabel metal2 32872 45640 32872 45640 0 _0273_
rlabel metal2 34664 45640 34664 45640 0 _0274_
rlabel metal2 45080 46368 45080 46368 0 _0275_
rlabel metal2 46984 46984 46984 46984 0 _0276_
rlabel metal2 49560 46200 49560 46200 0 _0277_
rlabel metal3 52080 45864 52080 45864 0 _0278_
rlabel metal2 50904 44688 50904 44688 0 _0279_
rlabel metal2 51072 43848 51072 43848 0 _0280_
rlabel metal2 9632 37240 9632 37240 0 _0281_
rlabel metal2 51240 43400 51240 43400 0 _0282_
rlabel metal2 50680 42952 50680 42952 0 _0283_
rlabel metal2 52696 43736 52696 43736 0 _0284_
rlabel metal2 39144 47656 39144 47656 0 _0285_
rlabel metal2 39536 49784 39536 49784 0 _0286_
rlabel metal2 30800 51912 30800 51912 0 _0287_
rlabel metal2 22456 54544 22456 54544 0 _0288_
rlabel metal4 22344 52192 22344 52192 0 _0289_
rlabel metal2 15176 51016 15176 51016 0 _0290_
rlabel metal2 12488 43064 12488 43064 0 _0291_
rlabel metal2 15680 47432 15680 47432 0 _0292_
rlabel metal2 15512 51296 15512 51296 0 _0293_
rlabel metal3 19208 50344 19208 50344 0 _0294_
rlabel metal2 22680 51016 22680 51016 0 _0295_
rlabel metal3 23128 47208 23128 47208 0 _0296_
rlabel metal2 24024 47488 24024 47488 0 _0297_
rlabel metal2 23464 47096 23464 47096 0 _0298_
rlabel metal3 39312 49112 39312 49112 0 _0299_
rlabel metal2 43960 48384 43960 48384 0 _0300_
rlabel metal2 51016 48608 51016 48608 0 _0301_
rlabel metal2 12376 45472 12376 45472 0 _0302_
rlabel metal2 33544 53592 33544 53592 0 _0303_
rlabel metal2 33320 52920 33320 52920 0 _0304_
rlabel metal2 32984 54488 32984 54488 0 _0305_
rlabel metal2 28056 54880 28056 54880 0 _0306_
rlabel metal2 16632 53424 16632 53424 0 _0307_
rlabel metal2 15848 52472 15848 52472 0 _0308_
rlabel metal2 19096 52584 19096 52584 0 _0309_
rlabel metal2 17024 52920 17024 52920 0 _0310_
rlabel metal3 30520 51352 30520 51352 0 _0311_
rlabel metal3 32648 51240 32648 51240 0 _0312_
rlabel metal2 31864 32872 31864 32872 0 _0313_
rlabel metal3 36232 51128 36232 51128 0 _0314_
rlabel metal3 46648 49784 46648 49784 0 _0315_
rlabel metal3 20440 47544 20440 47544 0 _0316_
rlabel metal2 29736 54880 29736 54880 0 _0317_
rlabel metal2 22288 54488 22288 54488 0 _0318_
rlabel metal2 30072 52136 30072 52136 0 _0319_
rlabel metal2 21504 49784 21504 49784 0 _0320_
rlabel metal3 36792 50008 36792 50008 0 _0321_
rlabel metal2 36456 49000 36456 49000 0 _0322_
rlabel metal2 35448 49616 35448 49616 0 _0323_
rlabel metal2 40040 34048 40040 34048 0 _0324_
rlabel metal2 50120 49392 50120 49392 0 _0325_
rlabel metal2 49784 48720 49784 48720 0 _0326_
rlabel metal2 50680 47768 50680 47768 0 _0327_
rlabel metal2 46144 45864 46144 45864 0 _0328_
rlabel metal2 47096 46144 47096 46144 0 _0329_
rlabel metal2 50456 47488 50456 47488 0 _0330_
rlabel metal2 51352 46984 51352 46984 0 _0331_
rlabel metal2 51352 45528 51352 45528 0 _0332_
rlabel metal2 51688 46312 51688 46312 0 _0333_
rlabel metal2 52920 46256 52920 46256 0 _0334_
rlabel metal2 51128 50960 51128 50960 0 _0335_
rlabel metal3 50008 48888 50008 48888 0 _0336_
rlabel metal2 50848 50456 50848 50456 0 _0337_
rlabel metal3 42224 46648 42224 46648 0 _0338_
rlabel metal2 43008 46760 43008 46760 0 _0339_
rlabel metal2 41160 51408 41160 51408 0 _0340_
rlabel metal2 27832 53592 27832 53592 0 _0341_
rlabel metal2 29288 50960 29288 50960 0 _0342_
rlabel metal3 25480 52136 25480 52136 0 _0343_
rlabel metal2 8568 10752 8568 10752 0 _0344_
rlabel metal2 28392 51408 28392 51408 0 _0345_
rlabel metal2 28000 51352 28000 51352 0 _0346_
rlabel metal2 27496 33516 27496 33516 0 _0347_
rlabel metal3 27944 50680 27944 50680 0 _0348_
rlabel metal2 27608 50456 27608 50456 0 _0349_
rlabel metal2 23128 52864 23128 52864 0 _0350_
rlabel metal2 27720 52080 27720 52080 0 _0351_
rlabel metal2 37576 51688 37576 51688 0 _0352_
rlabel metal2 38360 51072 38360 51072 0 _0353_
rlabel metal2 38808 50848 38808 50848 0 _0354_
rlabel metal2 10696 7952 10696 7952 0 _0355_
rlabel metal2 39256 50904 39256 50904 0 _0356_
rlabel metal2 42168 51240 42168 51240 0 _0357_
rlabel metal2 42504 50848 42504 50848 0 _0358_
rlabel metal2 23912 50904 23912 50904 0 _0359_
rlabel metal2 25368 51072 25368 51072 0 _0360_
rlabel metal3 22960 48104 22960 48104 0 _0361_
rlabel metal3 31920 51464 31920 51464 0 _0362_
rlabel metal2 42056 51408 42056 51408 0 _0363_
rlabel metal2 31752 51632 31752 51632 0 _0364_
rlabel metal2 26936 55692 26936 55692 0 _0365_
rlabel metal2 10696 14280 10696 14280 0 _0366_
rlabel metal2 19600 53032 19600 53032 0 _0367_
rlabel metal2 31976 53312 31976 53312 0 _0368_
rlabel metal2 34104 52472 34104 52472 0 _0369_
rlabel metal2 37240 54880 37240 54880 0 _0370_
rlabel metal2 34216 52584 34216 52584 0 _0371_
rlabel metal3 38696 52136 38696 52136 0 _0372_
rlabel metal2 43288 51744 43288 51744 0 _0373_
rlabel metal2 50456 50904 50456 50904 0 _0374_
rlabel metal2 51800 52584 51800 52584 0 _0375_
rlabel metal3 52360 50456 52360 50456 0 _0376_
rlabel metal2 5992 19152 5992 19152 0 _0377_
rlabel metal3 52304 50568 52304 50568 0 _0378_
rlabel metal2 52808 51072 52808 51072 0 _0379_
rlabel metal2 49896 46928 49896 46928 0 _0380_
rlabel metal3 51464 52080 51464 52080 0 _0381_
rlabel metal2 53424 51352 53424 51352 0 _0382_
rlabel metal3 38864 51352 38864 51352 0 _0383_
rlabel metal3 21392 52136 21392 52136 0 _0384_
rlabel metal2 22120 53592 22120 53592 0 _0385_
rlabel metal2 18984 49728 18984 49728 0 _0386_
rlabel metal2 6328 22008 6328 22008 0 _0387_
rlabel metal2 19320 50624 19320 50624 0 _0388_
rlabel metal2 22680 52472 22680 52472 0 _0389_
rlabel metal3 32088 52808 32088 52808 0 _0390_
rlabel metal3 40152 51912 40152 51912 0 _0391_
rlabel metal2 41608 52864 41608 52864 0 _0392_
rlabel metal2 31192 51856 31192 51856 0 _0393_
rlabel metal2 33320 48888 33320 48888 0 _0394_
rlabel metal2 35672 48608 35672 48608 0 _0395_
rlabel metal2 35784 49392 35784 49392 0 _0396_
rlabel metal2 37240 53648 37240 53648 0 _0397_
rlabel metal2 13888 16296 13888 16296 0 _0398_
rlabel metal2 34216 54096 34216 54096 0 _0399_
rlabel metal2 25480 52248 25480 52248 0 _0400_
rlabel metal2 26376 54824 26376 54824 0 _0401_
rlabel metal3 26432 53480 26432 53480 0 _0402_
rlabel metal3 24248 54488 24248 54488 0 _0403_
rlabel metal2 25816 53760 25816 53760 0 _0404_
rlabel metal2 26320 53704 26320 53704 0 _0405_
rlabel metal2 26824 54768 26824 54768 0 _0406_
rlabel metal2 27272 54488 27272 54488 0 _0407_
rlabel metal2 33040 55440 33040 55440 0 _0408_
rlabel metal2 12432 23352 12432 23352 0 _0409_
rlabel metal2 34776 54600 34776 54600 0 _0410_
rlabel metal2 36120 53760 36120 53760 0 _0411_
rlabel metal3 39704 53816 39704 53816 0 _0412_
rlabel metal2 43736 54040 43736 54040 0 _0413_
rlabel metal2 43848 54096 43848 54096 0 _0414_
rlabel metal2 49336 54544 49336 54544 0 _0415_
rlabel metal2 51352 53032 51352 53032 0 _0416_
rlabel metal3 52192 53592 52192 53592 0 _0417_
rlabel metal2 42056 53592 42056 53592 0 _0418_
rlabel metal2 12376 18536 12376 18536 0 _0419_
rlabel metal2 42280 54040 42280 54040 0 _0420_
rlabel metal2 24808 53984 24808 53984 0 _0421_
rlabel metal2 25144 53312 25144 53312 0 _0422_
rlabel metal2 31304 52696 31304 52696 0 _0423_
rlabel metal3 31444 52808 31444 52808 0 _0424_
rlabel metal2 39536 51576 39536 51576 0 _0425_
rlabel metal2 39032 54208 39032 54208 0 _0426_
rlabel metal2 34216 49000 34216 49000 0 _0427_
rlabel metal2 34496 50568 34496 50568 0 _0428_
rlabel metal3 32424 50456 32424 50456 0 _0429_
rlabel metal2 7784 15568 7784 15568 0 _0430_
rlabel metal3 33656 50568 33656 50568 0 _0431_
rlabel metal2 38136 53424 38136 53424 0 _0432_
rlabel metal2 28784 54488 28784 54488 0 _0433_
rlabel metal2 30968 53760 30968 53760 0 _0434_
rlabel metal2 31528 54320 31528 54320 0 _0435_
rlabel metal3 35560 55272 35560 55272 0 _0436_
rlabel metal2 39928 54488 39928 54488 0 _0437_
rlabel metal3 41776 55160 41776 55160 0 _0438_
rlabel metal2 44744 54712 44744 54712 0 _0439_
rlabel metal3 45192 55160 45192 55160 0 _0440_
rlabel metal3 10976 15400 10976 15400 0 _0441_
rlabel metal2 49112 54824 49112 54824 0 _0442_
rlabel metal3 46816 53592 46816 53592 0 _0443_
rlabel metal2 50232 54096 50232 54096 0 _0444_
rlabel metal2 51632 55272 51632 55272 0 _0445_
rlabel metal2 49224 53704 49224 53704 0 _0446_
rlabel metal2 47544 54320 47544 54320 0 _0447_
rlabel metal2 45192 54712 45192 54712 0 _0448_
rlabel metal3 46424 55160 46424 55160 0 _0449_
rlabel metal2 45192 50512 45192 50512 0 _0450_
rlabel metal2 18872 17752 18872 17752 0 _0451_
rlabel metal2 30632 54768 30632 54768 0 _0452_
rlabel metal2 34104 54432 34104 54432 0 _0453_
rlabel metal2 35616 55048 35616 55048 0 _0454_
rlabel metal2 44016 50568 44016 50568 0 _0455_
rlabel metal2 45808 51352 45808 51352 0 _0456_
rlabel metal2 29624 50176 29624 50176 0 _0457_
rlabel metal3 42280 49112 42280 49112 0 _0458_
rlabel metal2 42168 46928 42168 46928 0 _0459_
rlabel metal3 43064 49000 43064 49000 0 _0460_
rlabel metal3 43456 48888 43456 48888 0 _0461_
rlabel metal2 11144 21392 11144 21392 0 _0462_
rlabel metal2 45528 51072 45528 51072 0 _0463_
rlabel metal2 46424 52472 46424 52472 0 _0464_
rlabel metal2 38752 53032 38752 53032 0 _0465_
rlabel metal2 38920 53200 38920 53200 0 _0466_
rlabel metal2 46200 54152 46200 54152 0 _0467_
rlabel metal2 46872 54880 46872 54880 0 _0468_
rlabel metal2 47432 54768 47432 54768 0 _0469_
rlabel metal2 47712 55160 47712 55160 0 _0470_
rlabel metal2 46648 50512 46648 50512 0 _0471_
rlabel metal2 6272 20552 6272 20552 0 _0472_
rlabel metal3 46760 51464 46760 51464 0 _0473_
rlabel metal2 29904 51240 29904 51240 0 _0474_
rlabel metal2 39368 47264 39368 47264 0 _0475_
rlabel metal2 39760 47656 39760 47656 0 _0476_
rlabel metal2 40152 47600 40152 47600 0 _0477_
rlabel metal2 46032 49000 46032 49000 0 _0478_
rlabel metal2 46984 50904 46984 50904 0 _0479_
rlabel metal2 47880 52360 47880 52360 0 _0480_
rlabel metal2 47432 50848 47432 50848 0 _0481_
rlabel metal2 47992 53032 47992 53032 0 _0482_
rlabel metal2 6832 20552 6832 20552 0 _0483_
rlabel metal2 46984 53760 46984 53760 0 _0484_
rlabel metal2 47880 53760 47880 53760 0 _0485_
rlabel metal2 48944 53592 48944 53592 0 _0486_
rlabel metal2 48104 51576 48104 51576 0 _0487_
rlabel metal2 47768 49000 47768 49000 0 _0488_
rlabel metal2 46200 49280 46200 49280 0 _0489_
rlabel metal2 47544 48832 47544 48832 0 _0490_
rlabel metal2 47656 50568 47656 50568 0 _0491_
rlabel metal3 48328 50568 48328 50568 0 _0492_
rlabel metal3 9352 22344 9352 22344 0 _0493_
rlabel metal2 46536 36008 46536 36008 0 _0494_
rlabel metal2 43064 28504 43064 28504 0 _0495_
rlabel via1 23240 28392 23240 28392 0 _0496_
rlabel metal2 18424 28840 18424 28840 0 _0497_
rlabel metal2 12712 28952 12712 28952 0 _0498_
rlabel metal2 22960 26488 22960 26488 0 _0499_
rlabel metal2 12992 20776 12992 20776 0 _0500_
rlabel metal3 18704 27944 18704 27944 0 _0501_
rlabel metal3 18536 30072 18536 30072 0 _0502_
rlabel metal2 18760 30856 18760 30856 0 _0503_
rlabel metal2 24304 30968 24304 30968 0 _0504_
rlabel metal2 20440 29344 20440 29344 0 _0505_
rlabel metal3 25928 29960 25928 29960 0 _0506_
rlabel metal3 25032 30856 25032 30856 0 _0507_
rlabel metal2 10528 19880 10528 19880 0 _0508_
rlabel metal2 24024 31080 24024 31080 0 _0509_
rlabel metal2 23576 31416 23576 31416 0 _0510_
rlabel metal2 25368 30520 25368 30520 0 _0511_
rlabel metal2 26432 30408 26432 30408 0 _0512_
rlabel metal3 16492 25480 16492 25480 0 _0513_
rlabel metal2 18704 27944 18704 27944 0 _0514_
rlabel metal2 16744 23184 16744 23184 0 _0515_
rlabel metal2 20440 25872 20440 25872 0 _0516_
rlabel metal2 19656 25872 19656 25872 0 _0517_
rlabel metal2 25368 25760 25368 25760 0 _0518_
rlabel metal3 15624 26376 15624 26376 0 _0519_
rlabel metal2 23128 25872 23128 25872 0 _0520_
rlabel metal2 23744 26824 23744 26824 0 _0521_
rlabel metal2 24360 26544 24360 26544 0 _0522_
rlabel metal2 22904 25928 22904 25928 0 _0523_
rlabel metal2 14000 23912 14000 23912 0 _0524_
rlabel metal3 19432 25704 19432 25704 0 _0525_
rlabel metal2 22568 26628 22568 26628 0 _0526_
rlabel metal2 43120 33320 43120 33320 0 _0527_
rlabel metal2 14616 23464 14616 23464 0 _0528_
rlabel metal3 15736 25368 15736 25368 0 _0529_
rlabel metal2 15960 24360 15960 24360 0 _0530_
rlabel metal2 15288 24640 15288 24640 0 _0531_
rlabel metal2 16296 24248 16296 24248 0 _0532_
rlabel metal2 6776 19208 6776 19208 0 _0533_
rlabel metal2 6104 15792 6104 15792 0 _0534_
rlabel metal3 6720 12936 6720 12936 0 _0535_
rlabel metal3 8568 18424 8568 18424 0 _0536_
rlabel metal3 24360 20832 24360 20832 0 _0537_
rlabel metal2 15400 22848 15400 22848 0 _0538_
rlabel metal2 18648 23744 18648 23744 0 _0539_
rlabel metal2 22904 24360 22904 24360 0 _0540_
rlabel metal2 41496 16912 41496 16912 0 _0541_
rlabel metal2 30912 27832 30912 27832 0 _0542_
rlabel metal3 35168 30184 35168 30184 0 _0543_
rlabel metal3 36624 30296 36624 30296 0 _0544_
rlabel metal2 36232 41664 36232 41664 0 _0545_
rlabel metal2 35560 48664 35560 48664 0 _0546_
rlabel metal2 34104 27720 34104 27720 0 _0547_
rlabel metal2 39256 42728 39256 42728 0 _0548_
rlabel metal3 39480 50456 39480 50456 0 _0549_
rlabel metal2 31640 31360 31640 31360 0 _0550_
rlabel metal3 39256 26488 39256 26488 0 _0551_
rlabel metal2 37072 37352 37072 37352 0 _0552_
rlabel metal2 39480 33376 39480 33376 0 _0553_
rlabel metal3 38752 32536 38752 32536 0 _0554_
rlabel metal2 37912 32480 37912 32480 0 _0555_
rlabel metal2 40040 13888 40040 13888 0 _0556_
rlabel metal2 39592 20888 39592 20888 0 _0557_
rlabel metal3 39032 25368 39032 25368 0 _0558_
rlabel metal2 37912 26096 37912 26096 0 _0559_
rlabel metal2 39424 26264 39424 26264 0 _0560_
rlabel metal2 39368 26040 39368 26040 0 _0561_
rlabel metal2 39424 27832 39424 27832 0 _0562_
rlabel metal2 27776 28056 27776 28056 0 _0563_
rlabel metal2 29624 28672 29624 28672 0 _0564_
rlabel metal2 39144 29792 39144 29792 0 _0565_
rlabel metal2 44800 20552 44800 20552 0 _0566_
rlabel metal2 45416 19040 45416 19040 0 _0567_
rlabel metal2 17192 3920 17192 3920 0 _0568_
rlabel metal2 24472 5040 24472 5040 0 _0569_
rlabel metal2 26488 4592 26488 4592 0 _0570_
rlabel metal3 25200 16744 25200 16744 0 _0571_
rlabel metal2 7784 19992 7784 19992 0 _0572_
rlabel metal2 10808 16240 10808 16240 0 _0573_
rlabel metal3 16352 16296 16352 16296 0 _0574_
rlabel metal3 29232 15400 29232 15400 0 _0575_
rlabel metal3 6552 9240 6552 9240 0 _0576_
rlabel metal3 8092 3304 8092 3304 0 _0577_
rlabel metal2 26488 9800 26488 9800 0 _0578_
rlabel metal2 24248 6440 24248 6440 0 _0579_
rlabel metal3 28280 9240 28280 9240 0 _0580_
rlabel metal2 18312 19208 18312 19208 0 _0581_
rlabel metal2 16856 7616 16856 7616 0 _0582_
rlabel metal2 28616 9856 28616 9856 0 _0583_
rlabel metal2 8568 13216 8568 13216 0 _0584_
rlabel metal2 17864 19880 17864 19880 0 _0585_
rlabel metal2 13104 18536 13104 18536 0 _0586_
rlabel metal2 24472 14448 24472 14448 0 _0587_
rlabel metal2 26152 13104 26152 13104 0 _0588_
rlabel metal2 10248 12992 10248 12992 0 _0589_
rlabel metal3 14952 3304 14952 3304 0 _0590_
rlabel metal2 17864 17192 17864 17192 0 _0591_
rlabel metal2 19320 22064 19320 22064 0 _0592_
rlabel metal3 26432 20552 26432 20552 0 _0593_
rlabel metal2 29624 9520 29624 9520 0 _0594_
rlabel metal2 7504 10584 7504 10584 0 _0595_
rlabel metal3 17080 2744 17080 2744 0 _0596_
rlabel metal2 7336 17640 7336 17640 0 _0597_
rlabel metal2 9576 14560 9576 14560 0 _0598_
rlabel metal2 17584 7672 17584 7672 0 _0599_
rlabel metal2 24920 9464 24920 9464 0 _0600_
rlabel metal2 11480 16716 11480 16716 0 _0601_
rlabel metal3 23352 24192 23352 24192 0 _0602_
rlabel metal2 21448 6552 21448 6552 0 _0603_
rlabel metal2 10024 20048 10024 20048 0 _0604_
rlabel metal2 21784 18704 21784 18704 0 _0605_
rlabel metal2 25704 14224 25704 14224 0 _0606_
rlabel metal2 28056 23464 28056 23464 0 _0607_
rlabel metal2 29960 10472 29960 10472 0 _0608_
rlabel metal2 21448 12600 21448 12600 0 _0609_
rlabel metal3 27608 14280 27608 14280 0 _0610_
rlabel metal2 33096 17360 33096 17360 0 _0611_
rlabel metal2 15512 18312 15512 18312 0 _0612_
rlabel metal2 18760 19376 18760 19376 0 _0613_
rlabel metal2 24584 20552 24584 20552 0 _0614_
rlabel metal3 14504 3080 14504 3080 0 _0615_
rlabel metal2 25256 17304 25256 17304 0 _0616_
rlabel metal2 30520 18144 30520 18144 0 _0617_
rlabel metal2 39592 9912 39592 9912 0 _0618_
rlabel metal2 41272 5656 41272 5656 0 _0619_
rlabel metal3 16576 21560 16576 21560 0 _0620_
rlabel metal2 25536 24584 25536 24584 0 _0621_
rlabel metal2 33096 28952 33096 28952 0 _0622_
rlabel metal2 22008 17976 22008 17976 0 _0623_
rlabel metal3 7168 10584 7168 10584 0 _0624_
rlabel metal2 11816 7056 11816 7056 0 _0625_
rlabel metal2 10248 5488 10248 5488 0 _0626_
rlabel metal3 21896 5208 21896 5208 0 _0627_
rlabel metal2 26264 5208 26264 5208 0 _0628_
rlabel metal2 21112 8736 21112 8736 0 _0629_
rlabel metal2 12040 13440 12040 13440 0 _0630_
rlabel metal2 15288 8708 15288 8708 0 _0631_
rlabel metal2 14504 8008 14504 8008 0 _0632_
rlabel metal3 16968 15624 16968 15624 0 _0633_
rlabel metal3 19824 5096 19824 5096 0 _0634_
rlabel metal2 14168 6608 14168 6608 0 _0635_
rlabel metal2 15512 7504 15512 7504 0 _0636_
rlabel metal3 10416 5096 10416 5096 0 _0637_
rlabel metal2 14392 9744 14392 9744 0 _0638_
rlabel metal2 13160 9296 13160 9296 0 _0639_
rlabel metal2 17192 9408 17192 9408 0 _0640_
rlabel metal3 19712 24920 19712 24920 0 _0641_
rlabel metal2 24696 10528 24696 10528 0 _0642_
rlabel metal2 9352 22736 9352 22736 0 _0643_
rlabel metal2 17304 7616 17304 7616 0 _0644_
rlabel metal2 17976 7952 17976 7952 0 _0645_
rlabel metal2 17752 8960 17752 8960 0 _0646_
rlabel metal2 14504 14056 14504 14056 0 _0647_
rlabel metal2 7896 11368 7896 11368 0 _0648_
rlabel metal3 9576 15288 9576 15288 0 _0649_
rlabel metal2 14728 14392 14728 14392 0 _0650_
rlabel metal2 19600 10360 19600 10360 0 _0651_
rlabel metal2 15512 13720 15512 13720 0 _0652_
rlabel metal3 22008 3248 22008 3248 0 _0653_
rlabel metal3 43512 16072 43512 16072 0 _0654_
rlabel metal3 45192 16072 45192 16072 0 _0655_
rlabel metal2 47432 22512 47432 22512 0 _0656_
rlabel metal2 40264 6272 40264 6272 0 _0657_
rlabel metal2 39984 5880 39984 5880 0 _0658_
rlabel metal2 16184 18368 16184 18368 0 _0659_
rlabel metal2 21896 8960 21896 8960 0 _0660_
rlabel metal2 3304 15008 3304 15008 0 _0661_
rlabel metal2 24136 19936 24136 19936 0 _0662_
rlabel metal2 20776 20328 20776 20328 0 _0663_
rlabel metal2 15736 17416 15736 17416 0 _0664_
rlabel metal3 16912 15064 16912 15064 0 _0665_
rlabel metal3 23968 15960 23968 15960 0 _0666_
rlabel metal2 13384 16800 13384 16800 0 _0667_
rlabel metal2 16184 16688 16184 16688 0 _0668_
rlabel metal2 18872 19320 18872 19320 0 _0669_
rlabel metal2 21224 19264 21224 19264 0 _0670_
rlabel metal2 20104 19264 20104 19264 0 _0671_
rlabel metal2 10248 14616 10248 14616 0 _0672_
rlabel metal2 21672 17752 21672 17752 0 _0673_
rlabel metal2 19768 19712 19768 19712 0 _0674_
rlabel metal2 16296 19768 16296 19768 0 _0675_
rlabel metal2 19320 23968 19320 23968 0 _0676_
rlabel metal2 21448 23688 21448 23688 0 _0677_
rlabel metal2 19544 21560 19544 21560 0 _0678_
rlabel metal2 21112 23744 21112 23744 0 _0679_
rlabel metal2 38920 5432 38920 5432 0 _0680_
rlabel metal3 40264 5096 40264 5096 0 _0681_
rlabel metal3 40768 4312 40768 4312 0 _0682_
rlabel metal2 40096 5096 40096 5096 0 _0683_
rlabel metal2 42840 5152 42840 5152 0 _0684_
rlabel metal3 12432 3192 12432 3192 0 _0685_
rlabel metal2 22456 3808 22456 3808 0 _0686_
rlabel metal2 23016 5376 23016 5376 0 _0687_
rlabel metal2 24584 6048 24584 6048 0 _0688_
rlabel metal2 24472 7168 24472 7168 0 _0689_
rlabel metal2 20664 6552 20664 6552 0 _0690_
rlabel metal4 19432 6496 19432 6496 0 _0691_
rlabel metal3 20216 22064 20216 22064 0 _0692_
rlabel metal2 19096 7784 19096 7784 0 _0693_
rlabel metal2 20216 6328 20216 6328 0 _0694_
rlabel metal2 16744 19040 16744 19040 0 _0695_
rlabel metal2 21336 5656 21336 5656 0 _0696_
rlabel metal2 18536 5152 18536 5152 0 _0697_
rlabel metal3 15960 8904 15960 8904 0 _0698_
rlabel metal3 13720 9800 13720 9800 0 _0699_
rlabel metal2 23912 9408 23912 9408 0 _0700_
rlabel metal3 17416 8792 17416 8792 0 _0701_
rlabel metal3 20888 8792 20888 8792 0 _0702_
rlabel metal2 23464 5936 23464 5936 0 _0703_
rlabel metal2 39536 9240 39536 9240 0 _0704_
rlabel metal2 37128 7056 37128 7056 0 _0705_
rlabel metal2 41104 7448 41104 7448 0 _0706_
rlabel metal2 42840 13888 42840 13888 0 _0707_
rlabel metal2 39368 17976 39368 17976 0 _0708_
rlabel metal2 19768 13384 19768 13384 0 _0709_
rlabel metal2 19880 13384 19880 13384 0 _0710_
rlabel metal2 21000 13216 21000 13216 0 _0711_
rlabel metal2 25144 19488 25144 19488 0 _0712_
rlabel metal2 20104 22568 20104 22568 0 _0713_
rlabel metal2 19432 11984 19432 11984 0 _0714_
rlabel metal2 19208 11760 19208 11760 0 _0715_
rlabel metal2 18200 14224 18200 14224 0 _0716_
rlabel metal3 20272 11816 20272 11816 0 _0717_
rlabel metal3 11480 15960 11480 15960 0 _0718_
rlabel metal3 20776 12040 20776 12040 0 _0719_
rlabel metal3 17920 16072 17920 16072 0 _0720_
rlabel metal2 21000 15708 21000 15708 0 _0721_
rlabel metal2 19544 12880 19544 12880 0 _0722_
rlabel metal2 20440 3220 20440 3220 0 _0723_
rlabel metal2 40152 12544 40152 12544 0 _0724_
rlabel metal2 17192 19656 17192 19656 0 _0725_
rlabel metal2 10696 19488 10696 19488 0 _0726_
rlabel metal2 15288 10472 15288 10472 0 _0727_
rlabel metal2 17416 20552 17416 20552 0 _0728_
rlabel metal3 23296 21560 23296 21560 0 _0729_
rlabel metal2 14056 20552 14056 20552 0 _0730_
rlabel metal2 15848 13888 15848 13888 0 _0731_
rlabel metal3 14728 12936 14728 12936 0 _0732_
rlabel metal2 19768 15008 19768 15008 0 _0733_
rlabel metal3 26880 12600 26880 12600 0 _0734_
rlabel metal2 19208 3808 19208 3808 0 _0735_
rlabel metal2 13440 8232 13440 8232 0 _0736_
rlabel metal2 11592 12096 11592 12096 0 _0737_
rlabel metal2 17640 12656 17640 12656 0 _0738_
rlabel metal2 18312 12768 18312 12768 0 _0739_
rlabel metal2 14728 11032 14728 11032 0 _0740_
rlabel metal2 23352 12376 23352 12376 0 _0741_
rlabel metal2 17640 11088 17640 11088 0 _0742_
rlabel metal2 24136 21224 24136 21224 0 _0743_
rlabel metal2 16856 11592 16856 11592 0 _0744_
rlabel metal2 14616 8288 14616 8288 0 _0745_
rlabel metal3 8372 2856 8372 2856 0 _0746_
rlabel metal2 16408 9856 16408 9856 0 _0747_
rlabel metal2 25536 19992 25536 19992 0 _0748_
rlabel metal2 12824 9352 12824 9352 0 _0749_
rlabel metal2 15512 10080 15512 10080 0 _0750_
rlabel metal2 14952 9744 14952 9744 0 _0751_
rlabel metal4 18088 6328 18088 6328 0 _0752_
rlabel metal2 40040 12544 40040 12544 0 _0753_
rlabel metal2 41608 10192 41608 10192 0 _0754_
rlabel metal2 42616 6944 42616 6944 0 _0755_
rlabel metal3 42504 23240 42504 23240 0 _0756_
rlabel metal2 42840 21000 42840 21000 0 _0757_
rlabel metal2 41272 9688 41272 9688 0 _0758_
rlabel metal2 18200 18760 18200 18760 0 _0759_
rlabel via2 21448 4424 21448 4424 0 _0760_
rlabel metal2 24024 3976 24024 3976 0 _0761_
rlabel metal2 31416 20608 31416 20608 0 _0762_
rlabel metal2 9800 4760 9800 4760 0 _0763_
rlabel metal2 31976 7672 31976 7672 0 _0764_
rlabel metal2 26824 19656 26824 19656 0 _0765_
rlabel metal3 17752 16856 17752 16856 0 _0766_
rlabel metal2 30800 10472 30800 10472 0 _0767_
rlabel metal2 33600 8232 33600 8232 0 _0768_
rlabel metal2 30408 15400 30408 15400 0 _0769_
rlabel metal2 29064 7728 29064 7728 0 _0770_
rlabel metal2 30968 8680 30968 8680 0 _0771_
rlabel metal2 34328 10976 34328 10976 0 _0772_
rlabel metal2 34104 8680 34104 8680 0 _0773_
rlabel metal2 40600 9296 40600 9296 0 _0774_
rlabel metal2 42840 9408 42840 9408 0 _0775_
rlabel metal2 42840 7000 42840 7000 0 _0776_
rlabel metal3 45808 5096 45808 5096 0 _0777_
rlabel metal2 45528 5096 45528 5096 0 _0778_
rlabel metal2 40152 11032 40152 11032 0 _0779_
rlabel metal2 46760 6328 46760 6328 0 _0780_
rlabel metal2 19320 4592 19320 4592 0 _0781_
rlabel metal2 17976 4480 17976 4480 0 _0782_
rlabel metal2 17640 5096 17640 5096 0 _0783_
rlabel metal2 11368 2912 11368 2912 0 _0784_
rlabel metal3 17192 4536 17192 4536 0 _0785_
rlabel metal2 15400 5376 15400 5376 0 _0786_
rlabel metal2 14952 5152 14952 5152 0 _0787_
rlabel metal3 15960 5208 15960 5208 0 _0788_
rlabel metal2 17976 15568 17976 15568 0 _0789_
rlabel metal2 16072 6664 16072 6664 0 _0790_
rlabel metal3 16744 5320 16744 5320 0 _0791_
rlabel metal2 17752 2996 17752 2996 0 _0792_
rlabel metal2 37576 7896 37576 7896 0 _0793_
rlabel metal2 37912 7504 37912 7504 0 _0794_
rlabel metal2 43960 7392 43960 7392 0 _0795_
rlabel metal2 41384 16800 41384 16800 0 _0796_
rlabel metal2 45192 15904 45192 15904 0 _0797_
rlabel metal2 14056 16184 14056 16184 0 _0798_
rlabel metal2 14952 15232 14952 15232 0 _0799_
rlabel metal3 19264 13944 19264 13944 0 _0800_
rlabel metal2 18200 17192 18200 17192 0 _0801_
rlabel metal2 17640 16184 17640 16184 0 _0802_
rlabel metal3 19096 15064 19096 15064 0 _0803_
rlabel metal3 22512 15624 22512 15624 0 _0804_
rlabel metal2 18872 15904 18872 15904 0 _0805_
rlabel metal3 42280 15400 42280 15400 0 _0806_
rlabel metal3 42224 15288 42224 15288 0 _0807_
rlabel metal2 44632 9576 44632 9576 0 _0808_
rlabel metal2 44688 7448 44688 7448 0 _0809_
rlabel metal3 40264 8232 40264 8232 0 _0810_
rlabel metal2 20888 4928 20888 4928 0 _0811_
rlabel metal3 36960 20776 36960 20776 0 _0812_
rlabel metal2 31864 11648 31864 11648 0 _0813_
rlabel metal2 25760 3752 25760 3752 0 _0814_
rlabel metal3 32480 10696 32480 10696 0 _0815_
rlabel metal2 28504 7784 28504 7784 0 _0816_
rlabel metal2 25144 3920 25144 3920 0 _0817_
rlabel metal2 26600 17136 26600 17136 0 _0818_
rlabel metal3 31192 4200 31192 4200 0 _0819_
rlabel metal3 31584 5880 31584 5880 0 _0820_
rlabel metal2 30856 6216 30856 6216 0 _0821_
rlabel metal2 25480 18984 25480 18984 0 _0822_
rlabel metal3 22960 9912 22960 9912 0 _0823_
rlabel metal2 16072 9688 16072 9688 0 _0824_
rlabel metal3 22120 15288 22120 15288 0 _0825_
rlabel metal2 22960 3304 22960 3304 0 _0826_
rlabel metal3 26712 6552 26712 6552 0 _0827_
rlabel metal2 40376 7336 40376 7336 0 _0828_
rlabel metal2 41272 8568 41272 8568 0 _0829_
rlabel metal3 44912 7448 44912 7448 0 _0830_
rlabel metal2 46536 6048 46536 6048 0 _0831_
rlabel metal2 48384 5096 48384 5096 0 _0832_
rlabel metal2 46648 4928 46648 4928 0 _0833_
rlabel metal2 47544 5096 47544 5096 0 _0834_
rlabel metal2 50680 7112 50680 7112 0 _0835_
rlabel metal2 45864 7504 45864 7504 0 _0836_
rlabel metal2 45584 8120 45584 8120 0 _0837_
rlabel metal2 47992 6888 47992 6888 0 _0838_
rlabel metal2 26824 4928 26824 4928 0 _0839_
rlabel metal2 27888 11144 27888 11144 0 _0840_
rlabel metal2 28336 14280 28336 14280 0 _0841_
rlabel metal2 28952 12096 28952 12096 0 _0842_
rlabel metal2 29288 13216 29288 13216 0 _0843_
rlabel metal2 22568 13104 22568 13104 0 _0844_
rlabel metal2 23912 12824 23912 12824 0 _0845_
rlabel metal2 28280 8120 28280 8120 0 _0846_
rlabel metal2 21896 11648 21896 11648 0 _0847_
rlabel metal2 28280 12376 28280 12376 0 _0848_
rlabel metal2 25928 17752 25928 17752 0 _0849_
rlabel metal2 30408 12600 30408 12600 0 _0850_
rlabel metal2 35672 12600 35672 12600 0 _0851_
rlabel metal2 41272 12376 41272 12376 0 _0852_
rlabel metal2 22904 20944 22904 20944 0 _0853_
rlabel metal2 32088 5264 32088 5264 0 _0854_
rlabel metal2 33656 5880 33656 5880 0 _0855_
rlabel metal3 34608 7336 34608 7336 0 _0856_
rlabel metal2 42952 12096 42952 12096 0 _0857_
rlabel metal2 42952 10808 42952 10808 0 _0858_
rlabel metal2 42616 22008 42616 22008 0 _0859_
rlabel metal3 44128 10584 44128 10584 0 _0860_
rlabel metal2 43624 11144 43624 11144 0 _0861_
rlabel metal2 44856 10920 44856 10920 0 _0862_
rlabel metal2 47768 8288 47768 8288 0 _0863_
rlabel metal2 38248 19488 38248 19488 0 _0864_
rlabel metal2 37464 9072 37464 9072 0 _0865_
rlabel metal2 26096 18424 26096 18424 0 _0866_
rlabel metal2 24696 9968 24696 9968 0 _0867_
rlabel metal2 24248 11088 24248 11088 0 _0868_
rlabel metal2 27160 11648 27160 11648 0 _0869_
rlabel metal2 25312 20776 25312 20776 0 _0870_
rlabel metal2 25480 16296 25480 16296 0 _0871_
rlabel metal2 26040 11480 26040 11480 0 _0872_
rlabel metal2 26264 13328 26264 13328 0 _0873_
rlabel metal2 26712 23072 26712 23072 0 _0874_
rlabel metal2 26264 12488 26264 12488 0 _0875_
rlabel metal2 35896 10528 35896 10528 0 _0876_
rlabel metal2 46704 10584 46704 10584 0 _0877_
rlabel metal3 42672 13720 42672 13720 0 _0878_
rlabel metal2 21784 16240 21784 16240 0 _0879_
rlabel metal2 21616 14504 21616 14504 0 _0880_
rlabel metal2 21224 14616 21224 14616 0 _0881_
rlabel metal2 21784 6776 21784 6776 0 _0882_
rlabel metal2 24360 11648 24360 11648 0 _0883_
rlabel metal2 24472 11704 24472 11704 0 _0884_
rlabel metal3 21336 21672 21336 21672 0 _0885_
rlabel metal2 23520 11368 23520 11368 0 _0886_
rlabel metal2 36120 14056 36120 14056 0 _0887_
rlabel metal2 45528 14560 45528 14560 0 _0888_
rlabel metal2 46312 14448 46312 14448 0 _0889_
rlabel metal2 46648 13776 46648 13776 0 _0890_
rlabel metal2 47096 15904 47096 15904 0 _0891_
rlabel metal3 47824 17416 47824 17416 0 _0892_
rlabel metal2 47320 17360 47320 17360 0 _0893_
rlabel metal2 46984 15596 46984 15596 0 _0894_
rlabel metal2 48328 12992 48328 12992 0 _0895_
rlabel metal2 47880 8904 47880 8904 0 _0896_
rlabel metal2 46648 16772 46648 16772 0 _0897_
rlabel metal2 48440 10248 48440 10248 0 _0898_
rlabel metal2 49448 7840 49448 7840 0 _0899_
rlabel metal2 50568 7112 50568 7112 0 _0900_
rlabel metal2 51520 6552 51520 6552 0 _0901_
rlabel metal2 41944 11368 41944 11368 0 _0902_
rlabel metal2 29176 16912 29176 16912 0 _0903_
rlabel metal2 31976 13496 31976 13496 0 _0904_
rlabel metal2 30072 24080 30072 24080 0 _0905_
rlabel metal3 25144 23688 25144 23688 0 _0906_
rlabel metal3 19880 17528 19880 17528 0 _0907_
rlabel metal2 25816 18928 25816 18928 0 _0908_
rlabel metal2 30296 18704 30296 18704 0 _0909_
rlabel metal2 29848 17472 29848 17472 0 _0910_
rlabel metal2 27944 16240 27944 16240 0 _0911_
rlabel metal3 24024 19432 24024 19432 0 _0912_
rlabel metal2 26152 26152 26152 26152 0 _0913_
rlabel metal2 30072 15680 30072 15680 0 _0914_
rlabel metal2 31416 16576 31416 16576 0 _0915_
rlabel metal2 40376 15708 40376 15708 0 _0916_
rlabel metal2 43848 12488 43848 12488 0 _0917_
rlabel metal3 47768 12264 47768 12264 0 _0918_
rlabel metal2 38248 9800 38248 9800 0 _0919_
rlabel metal2 37576 11760 37576 11760 0 _0920_
rlabel metal2 28168 6552 28168 6552 0 _0921_
rlabel metal2 27216 5208 27216 5208 0 _0922_
rlabel metal3 26992 5208 26992 5208 0 _0923_
rlabel metal2 27720 5488 27720 5488 0 _0924_
rlabel metal2 31976 18032 31976 18032 0 _0925_
rlabel metal2 26320 19992 26320 19992 0 _0926_
rlabel metal2 32536 17920 32536 17920 0 _0927_
rlabel metal2 25816 13720 25816 13720 0 _0928_
rlabel metal2 33432 11256 33432 11256 0 _0929_
rlabel metal2 37688 10640 37688 10640 0 _0930_
rlabel metal2 46984 11760 46984 11760 0 _0931_
rlabel metal2 38136 16072 38136 16072 0 _0932_
rlabel metal2 38360 16128 38360 16128 0 _0933_
rlabel metal2 39144 16912 39144 16912 0 _0934_
rlabel metal2 38808 15932 38808 15932 0 _0935_
rlabel metal2 23912 22064 23912 22064 0 _0936_
rlabel metal2 33208 18536 33208 18536 0 _0937_
rlabel metal2 39704 19320 39704 19320 0 _0938_
rlabel metal2 33768 13384 33768 13384 0 _0939_
rlabel metal3 32928 17080 32928 17080 0 _0940_
rlabel metal2 23688 13160 23688 13160 0 _0941_
rlabel metal2 30856 12600 30856 12600 0 _0942_
rlabel metal2 32536 13776 32536 13776 0 _0943_
rlabel metal2 38696 14112 38696 14112 0 _0944_
rlabel metal2 26376 16184 26376 16184 0 _0945_
rlabel metal3 24472 16856 24472 16856 0 _0946_
rlabel metal2 22792 16352 22792 16352 0 _0947_
rlabel metal2 25256 23184 25256 23184 0 _0948_
rlabel metal2 22008 19936 22008 19936 0 _0949_
rlabel metal2 22848 16856 22848 16856 0 _0950_
rlabel metal2 25032 16296 25032 16296 0 _0951_
rlabel metal2 26264 16856 26264 16856 0 _0952_
rlabel metal2 22568 17304 22568 17304 0 _0953_
rlabel metal2 39592 16464 39592 16464 0 _0954_
rlabel metal3 39816 14952 39816 14952 0 _0955_
rlabel metal2 47432 12320 47432 12320 0 _0956_
rlabel metal3 48496 11368 48496 11368 0 _0957_
rlabel metal3 48552 12152 48552 12152 0 _0958_
rlabel metal2 50568 10136 50568 10136 0 _0959_
rlabel metal2 51800 13384 51800 13384 0 _0960_
rlabel metal2 50456 11592 50456 11592 0 _0961_
rlabel metal2 47880 10528 47880 10528 0 _0962_
rlabel metal2 51016 10248 51016 10248 0 _0963_
rlabel metal2 51800 9800 51800 9800 0 _0964_
rlabel metal2 50232 10080 50232 10080 0 _0965_
rlabel metal2 52024 9296 52024 9296 0 _0966_
rlabel metal2 49000 7728 49000 7728 0 _0967_
rlabel metal2 48888 7728 48888 7728 0 _0968_
rlabel metal3 50400 7448 50400 7448 0 _0969_
rlabel metal2 52752 10472 52752 10472 0 _0970_
rlabel metal2 53536 9016 53536 9016 0 _0971_
rlabel metal2 51016 12544 51016 12544 0 _0972_
rlabel metal3 52192 12936 52192 12936 0 _0973_
rlabel metal3 27384 22456 27384 22456 0 _0974_
rlabel metal2 26152 4088 26152 4088 0 _0975_
rlabel metal2 28336 10024 28336 10024 0 _0976_
rlabel metal2 35672 10696 35672 10696 0 _0977_
rlabel metal2 32200 11256 32200 11256 0 _0978_
rlabel metal2 32424 11088 32424 11088 0 _0979_
rlabel metal2 36232 10920 36232 10920 0 _0980_
rlabel metal2 35896 12600 35896 12600 0 _0981_
rlabel metal3 37688 11480 37688 11480 0 _0982_
rlabel metal2 48888 15148 48888 15148 0 _0983_
rlabel metal2 39928 17360 39928 17360 0 _0984_
rlabel metal2 20888 10304 20888 10304 0 _0985_
rlabel metal2 24024 11088 24024 11088 0 _0986_
rlabel metal2 23632 17528 23632 17528 0 _0987_
rlabel metal2 19320 9520 19320 9520 0 _0988_
rlabel metal2 19544 8120 19544 8120 0 _0989_
rlabel metal3 19152 10472 19152 10472 0 _0990_
rlabel metal2 19992 8680 19992 8680 0 _0991_
rlabel metal2 20440 10304 20440 10304 0 _0992_
rlabel metal2 39032 17304 39032 17304 0 _0993_
rlabel metal2 37856 16296 37856 16296 0 _0994_
rlabel metal2 48216 16352 48216 16352 0 _0995_
rlabel metal3 47376 16072 47376 16072 0 _0996_
rlabel metal3 48608 15848 48608 15848 0 _0997_
rlabel metal2 40152 22568 40152 22568 0 _0998_
rlabel metal2 42280 18816 42280 18816 0 _0999_
rlabel metal2 41664 21336 41664 21336 0 _1000_
rlabel metal3 26320 22232 26320 22232 0 _1001_
rlabel metal3 30576 21784 30576 21784 0 _1002_
rlabel metal2 33768 20048 33768 20048 0 _1003_
rlabel metal2 34104 20384 34104 20384 0 _1004_
rlabel metal2 25816 21840 25816 21840 0 _1005_
rlabel metal3 25200 21448 25200 21448 0 _1006_
rlabel metal2 21000 24080 21000 24080 0 _1007_
rlabel metal2 23856 16968 23856 16968 0 _1008_
rlabel metal3 24192 21784 24192 21784 0 _1009_
rlabel metal2 26600 21112 26600 21112 0 _1010_
rlabel metal2 41608 20720 41608 20720 0 _1011_
rlabel metal2 41832 21784 41832 21784 0 _1012_
rlabel metal3 46032 16184 46032 16184 0 _1013_
rlabel metal2 52248 14112 52248 14112 0 _1014_
rlabel metal3 54264 12152 54264 12152 0 _1015_
rlabel metal2 52136 11480 52136 11480 0 _1016_
rlabel metal2 53200 10472 53200 10472 0 _1017_
rlabel metal2 53984 10472 53984 10472 0 _1018_
rlabel metal2 55440 12152 55440 12152 0 _1019_
rlabel metal2 42952 17808 42952 17808 0 _1020_
rlabel metal3 28112 19208 28112 19208 0 _1021_
rlabel metal2 29232 19208 29232 19208 0 _1022_
rlabel metal2 21672 19656 21672 19656 0 _1023_
rlabel metal3 17360 19992 17360 19992 0 _1024_
rlabel metal2 18088 19264 18088 19264 0 _1025_
rlabel metal3 19880 20104 19880 20104 0 _1026_
rlabel metal2 21784 20440 21784 20440 0 _1027_
rlabel metal2 43960 18872 43960 18872 0 _1028_
rlabel metal2 44856 18480 44856 18480 0 _1029_
rlabel metal3 48104 18424 48104 18424 0 _1030_
rlabel metal2 37912 19320 37912 19320 0 _1031_
rlabel metal2 37576 22232 37576 22232 0 _1032_
rlabel metal2 22008 22008 22008 22008 0 _1033_
rlabel metal2 21784 22064 21784 22064 0 _1034_
rlabel metal2 29736 21840 29736 21840 0 _1035_
rlabel metal2 30968 23520 30968 23520 0 _1036_
rlabel metal2 31080 22008 31080 22008 0 _1037_
rlabel metal3 34272 21336 34272 21336 0 _1038_
rlabel metal2 49224 19712 49224 19712 0 _1039_
rlabel metal2 51072 19208 51072 19208 0 _1040_
rlabel metal2 44184 21784 44184 21784 0 _1041_
rlabel metal3 44744 22120 44744 22120 0 _1042_
rlabel metal3 33432 21672 33432 21672 0 _1043_
rlabel metal2 31976 19264 31976 19264 0 _1044_
rlabel metal2 23856 23800 23856 23800 0 _1045_
rlabel metal2 28728 24920 28728 24920 0 _1046_
rlabel metal2 28560 23128 28560 23128 0 _1047_
rlabel metal2 25648 23240 25648 23240 0 _1048_
rlabel metal3 28056 23128 28056 23128 0 _1049_
rlabel metal2 30296 22624 30296 22624 0 _1050_
rlabel metal2 26544 24584 26544 24584 0 _1051_
rlabel metal2 30072 22680 30072 22680 0 _1052_
rlabel metal2 44520 22848 44520 22848 0 _1053_
rlabel metal2 44576 23352 44576 23352 0 _1054_
rlabel metal2 46200 21784 46200 21784 0 _1055_
rlabel metal3 52248 16072 52248 16072 0 _1056_
rlabel metal3 50232 15288 50232 15288 0 _1057_
rlabel metal2 51240 15680 51240 15680 0 _1058_
rlabel metal2 50344 15176 50344 15176 0 _1059_
rlabel metal3 52416 16184 52416 16184 0 _1060_
rlabel metal2 53592 15344 53592 15344 0 _1061_
rlabel metal2 52360 12432 52360 12432 0 _1062_
rlabel metal2 51912 12992 51912 12992 0 _1063_
rlabel metal2 53088 12264 53088 12264 0 _1064_
rlabel metal2 54264 14840 54264 14840 0 _1065_
rlabel metal2 36232 20776 36232 20776 0 _1066_
rlabel metal2 33320 24248 33320 24248 0 _1067_
rlabel metal2 31192 20496 31192 20496 0 _1068_
rlabel metal2 32312 21336 32312 21336 0 _1069_
rlabel metal2 32704 21784 32704 21784 0 _1070_
rlabel metal2 33096 22400 33096 22400 0 _1071_
rlabel metal2 36008 21672 36008 21672 0 _1072_
rlabel metal2 49448 21280 49448 21280 0 _1073_
rlabel metal2 41832 17864 41832 17864 0 _1074_
rlabel metal2 30184 25480 30184 25480 0 _1075_
rlabel metal2 34216 14448 34216 14448 0 _1076_
rlabel metal2 33880 14952 33880 14952 0 _1077_
rlabel metal3 29288 15736 29288 15736 0 _1078_
rlabel metal2 32200 15232 32200 15232 0 _1079_
rlabel metal2 34216 15400 34216 15400 0 _1080_
rlabel metal2 34664 16128 34664 16128 0 _1081_
rlabel metal2 34328 16296 34328 16296 0 _1082_
rlabel metal2 34776 16968 34776 16968 0 _1083_
rlabel metal2 40936 17136 40936 17136 0 _1084_
rlabel metal3 44520 17416 44520 17416 0 _1085_
rlabel metal2 43400 15680 43400 15680 0 _1086_
rlabel metal2 45528 16576 45528 16576 0 _1087_
rlabel metal2 46424 17192 46424 17192 0 _1088_
rlabel metal2 49672 20440 49672 20440 0 _1089_
rlabel metal2 38192 22232 38192 22232 0 _1090_
rlabel metal2 29848 25032 29848 25032 0 _1091_
rlabel metal2 30520 24192 30520 24192 0 _1092_
rlabel metal2 37800 23072 37800 23072 0 _1093_
rlabel metal2 43736 22400 43736 22400 0 _1094_
rlabel metal2 44072 21952 44072 21952 0 _1095_
rlabel metal3 47040 22344 47040 22344 0 _1096_
rlabel metal3 51408 18424 51408 18424 0 _1097_
rlabel metal2 49560 18144 49560 18144 0 _1098_
rlabel metal2 50904 18816 50904 18816 0 _1099_
rlabel metal2 53368 16800 53368 16800 0 _1100_
rlabel metal2 52136 17416 52136 17416 0 _1101_
rlabel metal2 52808 16072 52808 16072 0 _1102_
rlabel metal2 54376 17416 54376 17416 0 _1103_
rlabel metal2 55048 17192 55048 17192 0 _1104_
rlabel metal2 35168 19992 35168 19992 0 _1105_
rlabel metal2 37016 19768 37016 19768 0 _1106_
rlabel metal2 46648 20496 46648 20496 0 _1107_
rlabel metal2 34888 17640 34888 17640 0 _1108_
rlabel metal2 24696 12824 24696 12824 0 _1109_
rlabel metal2 23016 12992 23016 12992 0 _1110_
rlabel metal2 24136 16408 24136 16408 0 _1111_
rlabel metal2 25144 13216 25144 13216 0 _1112_
rlabel metal2 41048 18088 41048 18088 0 _1113_
rlabel metal2 42168 18704 42168 18704 0 _1114_
rlabel metal2 46424 20048 46424 20048 0 _1115_
rlabel metal2 47544 22064 47544 22064 0 _1116_
rlabel metal2 23016 26040 23016 26040 0 _1117_
rlabel metal2 39480 22120 39480 22120 0 _1118_
rlabel metal2 30856 25928 30856 25928 0 _1119_
rlabel metal2 39200 22568 39200 22568 0 _1120_
rlabel metal2 40152 20664 40152 20664 0 _1121_
rlabel metal2 39928 21504 39928 21504 0 _1122_
rlabel metal2 40040 22848 40040 22848 0 _1123_
rlabel metal3 40544 23128 40544 23128 0 _1124_
rlabel metal2 47320 22736 47320 22736 0 _1125_
rlabel metal3 47992 22624 47992 22624 0 _1126_
rlabel metal2 50568 21336 50568 21336 0 _1127_
rlabel metal2 50008 21448 50008 21448 0 _1128_
rlabel metal2 51016 21728 51016 21728 0 _1129_
rlabel metal2 53368 21168 53368 21168 0 _1130_
rlabel metal2 54320 21672 54320 21672 0 _1131_
rlabel metal2 53368 19208 53368 19208 0 _1132_
rlabel metal2 52584 18088 52584 18088 0 _1133_
rlabel metal2 53256 17808 53256 17808 0 _1134_
rlabel metal2 52248 11704 52248 11704 0 _1135_
rlabel metal2 54376 11704 54376 11704 0 _1136_
rlabel metal2 53760 18424 53760 18424 0 _1137_
rlabel metal2 54264 19656 54264 19656 0 _1138_
rlabel metal2 54656 20664 54656 20664 0 _1139_
rlabel metal2 47600 21000 47600 21000 0 _1140_
rlabel metal2 46872 21336 46872 21336 0 _1141_
rlabel metal2 47656 22512 47656 22512 0 _1142_
rlabel metal2 35672 23128 35672 23128 0 _1143_
rlabel metal2 35616 24136 35616 24136 0 _1144_
rlabel metal2 24808 25424 24808 25424 0 _1145_
rlabel metal2 34216 25480 34216 25480 0 _1146_
rlabel metal2 34552 24528 34552 24528 0 _1147_
rlabel metal2 35840 24472 35840 24472 0 _1148_
rlabel metal2 47992 23744 47992 23744 0 _1149_
rlabel metal3 25088 23912 25088 23912 0 _1150_
rlabel metal2 26096 23912 26096 23912 0 _1151_
rlabel metal2 28392 23744 28392 23744 0 _1152_
rlabel metal2 41608 20216 41608 20216 0 _1153_
rlabel metal2 41944 19488 41944 19488 0 _1154_
rlabel metal2 46984 19544 46984 19544 0 _1155_
rlabel metal2 48216 23968 48216 23968 0 _1156_
rlabel metal2 48888 24080 48888 24080 0 _1157_
rlabel metal2 49784 24192 49784 24192 0 _1158_
rlabel metal3 19208 23800 19208 23800 0 _1159_
rlabel metal2 33768 24696 33768 24696 0 _1160_
rlabel metal2 43176 24416 43176 24416 0 _1161_
rlabel metal2 43512 24416 43512 24416 0 _1162_
rlabel metal2 49336 24304 49336 24304 0 _1163_
rlabel metal2 50232 23576 50232 23576 0 _1164_
rlabel metal2 52752 23352 52752 23352 0 _1165_
rlabel metal2 52920 24304 52920 24304 0 _1166_
rlabel metal2 53256 24472 53256 24472 0 _1167_
rlabel metal2 53928 22400 53928 22400 0 _1168_
rlabel metal2 53592 21840 53592 21840 0 _1169_
rlabel metal2 53816 22512 53816 22512 0 _1170_
rlabel metal2 54544 23240 54544 23240 0 _1171_
rlabel metal2 36792 23632 36792 23632 0 _1172_
rlabel metal2 46536 25368 46536 25368 0 _1173_
rlabel metal2 34944 21784 34944 21784 0 _1174_
rlabel metal3 32928 23128 32928 23128 0 _1175_
rlabel metal2 45416 23240 45416 23240 0 _1176_
rlabel metal2 45640 21504 45640 21504 0 _1177_
rlabel metal2 44856 23520 44856 23520 0 _1178_
rlabel metal3 45752 25480 45752 25480 0 _1179_
rlabel metal2 49112 25928 49112 25928 0 _1180_
rlabel metal2 25816 25144 25816 25144 0 _1181_
rlabel metal2 42392 25536 42392 25536 0 _1182_
rlabel metal2 43064 25536 43064 25536 0 _1183_
rlabel metal2 42616 25984 42616 25984 0 _1184_
rlabel metal2 43512 26488 43512 26488 0 _1185_
rlabel metal2 46480 26824 46480 26824 0 _1186_
rlabel metal3 50064 26376 50064 26376 0 _1187_
rlabel metal2 49504 23352 49504 23352 0 _1188_
rlabel metal2 48888 25200 48888 25200 0 _1189_
rlabel metal2 51632 25592 51632 25592 0 _1190_
rlabel metal2 52976 26824 52976 26824 0 _1191_
rlabel metal2 53032 23688 53032 23688 0 _1192_
rlabel metal2 53592 26096 53592 26096 0 _1193_
rlabel metal2 54544 26264 54544 26264 0 _1194_
rlabel metal2 47152 26488 47152 26488 0 _1195_
rlabel metal2 49448 27552 49448 27552 0 _1196_
rlabel metal2 49728 27272 49728 27272 0 _1197_
rlabel metal2 34944 18424 34944 18424 0 _1198_
rlabel metal2 43288 18144 43288 18144 0 _1199_
rlabel via2 22232 33096 22232 33096 0 _1200_
rlabel metal2 43624 18536 43624 18536 0 _1201_
rlabel metal3 43960 17528 43960 17528 0 _1202_
rlabel metal2 45528 18144 45528 18144 0 _1203_
rlabel metal2 46704 26376 46704 26376 0 _1204_
rlabel metal3 48944 27720 48944 27720 0 _1205_
rlabel metal2 52024 26572 52024 26572 0 _1206_
rlabel metal3 51016 27608 51016 27608 0 _1207_
rlabel metal3 52472 27832 52472 27832 0 _1208_
rlabel metal2 50680 26264 50680 26264 0 _1209_
rlabel metal2 53144 27440 53144 27440 0 _1210_
rlabel metal2 14504 34048 14504 34048 0 _1211_
rlabel metal2 53760 27832 53760 27832 0 _1212_
rlabel metal2 46144 26376 46144 26376 0 _1213_
rlabel metal2 46312 26712 46312 26712 0 _1214_
rlabel metal2 45976 25480 45976 25480 0 _1215_
rlabel metal2 50120 26600 50120 26600 0 _1216_
rlabel metal3 51912 26264 51912 26264 0 _1217_
rlabel metal2 46984 24640 46984 24640 0 _1218_
rlabel metal2 43680 5096 43680 5096 0 _1219_
rlabel metal2 21448 40544 21448 40544 0 _1220_
rlabel metal2 14392 31192 14392 31192 0 _1221_
rlabel metal2 14952 34608 14952 34608 0 _1222_
rlabel metal3 16296 43624 16296 43624 0 _1223_
rlabel metal2 19432 35392 19432 35392 0 _1224_
rlabel metal2 18648 33320 18648 33320 0 _1225_
rlabel metal2 16856 40208 16856 40208 0 _1226_
rlabel metal2 32200 37576 32200 37576 0 _1227_
rlabel metal3 23016 33320 23016 33320 0 _1228_
rlabel metal3 21280 37016 21280 37016 0 _1229_
rlabel metal2 24136 49840 24136 49840 0 _1230_
rlabel metal2 22904 42112 22904 42112 0 _1231_
rlabel metal2 12152 32760 12152 32760 0 _1232_
rlabel metal2 18088 40712 18088 40712 0 _1233_
rlabel metal2 16856 34496 16856 34496 0 _1234_
rlabel metal2 16072 46928 16072 46928 0 _1235_
rlabel metal2 19208 41608 19208 41608 0 _1236_
rlabel metal2 16184 38920 16184 38920 0 _1237_
rlabel metal2 9856 39704 9856 39704 0 _1238_
rlabel metal2 13496 43232 13496 43232 0 _1239_
rlabel metal2 24248 40768 24248 40768 0 _1240_
rlabel metal3 9520 31752 9520 31752 0 _1241_
rlabel metal2 26040 42168 26040 42168 0 _1242_
rlabel metal3 24584 41608 24584 41608 0 _1243_
rlabel metal2 21560 40040 21560 40040 0 _1244_
rlabel metal3 10584 34216 10584 34216 0 _1245_
rlabel metal2 10864 33320 10864 33320 0 _1246_
rlabel metal3 9688 36344 9688 36344 0 _1247_
rlabel metal3 20776 40936 20776 40936 0 _1248_
rlabel metal2 15008 36456 15008 36456 0 _1249_
rlabel metal2 24864 40376 24864 40376 0 _1250_
rlabel metal2 7896 36512 7896 36512 0 _1251_
rlabel metal2 11480 31892 11480 31892 0 _1252_
rlabel metal3 12040 35784 12040 35784 0 _1253_
rlabel metal2 27608 36008 27608 36008 0 _1254_
rlabel metal2 22456 40320 22456 40320 0 _1255_
rlabel metal2 28056 45360 28056 45360 0 _1256_
rlabel metal2 29176 35784 29176 35784 0 _1257_
rlabel metal2 29848 37072 29848 37072 0 _1258_
rlabel metal2 29400 40936 29400 40936 0 _1259_
rlabel metal2 39032 40544 39032 40544 0 _1260_
rlabel metal2 14840 35056 14840 35056 0 _1261_
rlabel metal2 27104 36904 27104 36904 0 _1262_
rlabel metal2 11368 46648 11368 46648 0 _1263_
rlabel metal2 17976 50120 17976 50120 0 _1264_
rlabel metal2 13496 40936 13496 40936 0 _1265_
rlabel metal2 16856 41608 16856 41608 0 _1266_
rlabel metal2 19152 39592 19152 39592 0 _1267_
rlabel metal2 17752 39088 17752 39088 0 _1268_
rlabel metal2 18256 47208 18256 47208 0 _1269_
rlabel metal2 17528 43512 17528 43512 0 _1270_
rlabel metal2 19432 39816 19432 39816 0 _1271_
rlabel metal2 11200 33096 11200 33096 0 _1272_
rlabel metal2 27160 33544 27160 33544 0 _1273_
rlabel metal2 13496 50624 13496 50624 0 _1274_
rlabel metal2 28224 32984 28224 32984 0 _1275_
rlabel metal2 28448 36680 28448 36680 0 _1276_
rlabel metal2 39144 39984 39144 39984 0 _1277_
rlabel metal3 40768 40488 40768 40488 0 _1278_
rlabel metal3 42952 38808 42952 38808 0 _1279_
rlabel metal2 42280 39592 42280 39592 0 _1280_
rlabel metal2 43512 41552 43512 41552 0 _1281_
rlabel metal2 43960 38024 43960 38024 0 _1282_
rlabel metal2 32200 40880 32200 40880 0 _1283_
rlabel metal2 23800 37632 23800 37632 0 _1284_
rlabel metal2 12712 33712 12712 33712 0 _1285_
rlabel metal2 26376 37464 26376 37464 0 _1286_
rlabel metal3 20720 38920 20720 38920 0 _1287_
rlabel metal3 19208 33544 19208 33544 0 _1288_
rlabel metal2 29288 34944 29288 34944 0 _1289_
rlabel metal3 25424 38696 25424 38696 0 _1290_
rlabel metal2 26936 37800 26936 37800 0 _1291_
rlabel metal3 12432 31864 12432 31864 0 _1292_
rlabel metal2 23912 42336 23912 42336 0 _1293_
rlabel metal3 31304 39032 31304 39032 0 _1294_
rlabel metal3 13944 38024 13944 38024 0 _1295_
rlabel metal2 25592 36288 25592 36288 0 _1296_
rlabel metal2 31136 38136 31136 38136 0 _1297_
rlabel metal2 30632 38864 30632 38864 0 _1298_
rlabel metal3 31136 39592 31136 39592 0 _1299_
rlabel metal2 15512 41720 15512 41720 0 _1300_
rlabel metal3 22344 39704 22344 39704 0 _1301_
rlabel metal2 24136 32480 24136 32480 0 _1302_
rlabel metal2 24416 42280 24416 42280 0 _1303_
rlabel metal2 23912 38920 23912 38920 0 _1304_
rlabel metal2 31192 39536 31192 39536 0 _1305_
rlabel metal2 36904 37128 36904 37128 0 _1306_
rlabel metal2 11256 32704 11256 32704 0 _1307_
rlabel metal2 42056 36512 42056 36512 0 _1308_
rlabel metal2 26152 34048 26152 34048 0 _1309_
rlabel metal2 11704 33824 11704 33824 0 _1310_
rlabel metal2 26376 34384 26376 34384 0 _1311_
rlabel metal2 27048 34720 27048 34720 0 _1312_
rlabel metal2 28728 33992 28728 33992 0 _1313_
rlabel metal2 30072 34664 30072 34664 0 _1314_
rlabel metal2 27496 36512 27496 36512 0 _1315_
rlabel metal2 27832 55104 27832 55104 0 _1316_
rlabel metal2 33880 35784 33880 35784 0 _1317_
rlabel metal2 24360 37744 24360 37744 0 _1318_
rlabel metal2 34216 35952 34216 35952 0 _1319_
rlabel metal2 42448 36456 42448 36456 0 _1320_
rlabel metal2 43512 36008 43512 36008 0 _1321_
rlabel metal2 44520 36008 44520 36008 0 _1322_
rlabel metal2 31192 34272 31192 34272 0 _1323_
rlabel metal2 26040 44744 26040 44744 0 _1324_
rlabel metal2 17416 45360 17416 45360 0 _1325_
rlabel metal2 23016 43064 23016 43064 0 _1326_
rlabel metal2 19824 42728 19824 42728 0 _1327_
rlabel metal3 28728 37800 28728 37800 0 _1328_
rlabel metal2 16072 38752 16072 38752 0 _1329_
rlabel metal2 18424 43344 18424 43344 0 _1330_
rlabel metal2 19544 43904 19544 43904 0 _1331_
rlabel metal3 22680 43288 22680 43288 0 _1332_
rlabel metal2 27048 43288 27048 43288 0 _1333_
rlabel metal2 17136 42616 17136 42616 0 _1334_
rlabel metal2 18200 42784 18200 42784 0 _1335_
rlabel metal3 25816 45192 25816 45192 0 _1336_
rlabel metal3 23016 42728 23016 42728 0 _1337_
rlabel metal2 8344 36512 8344 36512 0 _1338_
rlabel metal2 27048 37128 27048 37128 0 _1339_
rlabel metal2 9016 37464 9016 37464 0 _1340_
rlabel metal3 25312 45080 25312 45080 0 _1341_
rlabel metal2 24472 44576 24472 44576 0 _1342_
rlabel metal2 25256 42448 25256 42448 0 _1343_
rlabel metal2 26600 45304 26600 45304 0 _1344_
rlabel metal3 13776 48216 13776 48216 0 _1345_
rlabel metal2 15512 49168 15512 49168 0 _1346_
rlabel metal2 28168 53368 28168 53368 0 _1347_
rlabel metal2 24192 46872 24192 46872 0 _1348_
rlabel metal2 25032 44576 25032 44576 0 _1349_
rlabel metal3 11144 31192 11144 31192 0 _1350_
rlabel metal3 19488 45864 19488 45864 0 _1351_
rlabel metal2 39256 43344 39256 43344 0 _1352_
rlabel metal2 40600 39480 40600 39480 0 _1353_
rlabel metal2 41384 39592 41384 39592 0 _1354_
rlabel metal2 41048 39004 41048 39004 0 _1355_
rlabel metal2 24136 33320 24136 33320 0 _1356_
rlabel metal2 24696 33488 24696 33488 0 _1357_
rlabel metal3 24976 40488 24976 40488 0 _1358_
rlabel metal2 15736 42336 15736 42336 0 _1359_
rlabel metal3 13440 38136 13440 38136 0 _1360_
rlabel metal2 11480 37408 11480 37408 0 _1361_
rlabel metal2 20440 40600 20440 40600 0 _1362_
rlabel metal2 25648 39592 25648 39592 0 _1363_
rlabel metal2 23688 42336 23688 42336 0 _1364_
rlabel metal2 25256 40880 25256 40880 0 _1365_
rlabel metal2 26264 40656 26264 40656 0 _1366_
rlabel metal3 26376 36288 26376 36288 0 _1367_
rlabel metal2 20328 40264 20328 40264 0 _1368_
rlabel metal2 29624 39872 29624 39872 0 _1369_
rlabel metal3 25144 38808 25144 38808 0 _1370_
rlabel metal2 27384 51408 27384 51408 0 _1371_
rlabel metal2 14840 29960 14840 29960 0 _1372_
rlabel metal3 1358 28952 1358 28952 0 addI[0]
rlabel metal3 1358 30968 1358 30968 0 addI[1]
rlabel metal3 1358 32984 1358 32984 0 addI[2]
rlabel metal3 1358 31640 1358 31640 0 addI[3]
rlabel metal3 1358 33656 1358 33656 0 addI[4]
rlabel metal2 29624 57610 29624 57610 0 addI[5]
rlabel metal3 1358 21560 1358 21560 0 addQ[0]
rlabel metal3 1358 22904 1358 22904 0 addQ[1]
rlabel metal3 1358 22232 1358 22232 0 addQ[2]
rlabel metal3 1358 23576 1358 23576 0 addQ[3]
rlabel metal3 1358 26264 1358 26264 0 addQ[4]
rlabel metal3 1358 24248 1358 24248 0 addQ[5]
rlabel metal2 30352 28616 30352 28616 0 gen_sym.Reg_2M.data_in
rlabel metal2 33320 30576 33320 30576 0 gen_sym.Reg_2M.data_out
rlabel metal2 29848 29904 29848 29904 0 gen_sym.Reg_2M.enable
rlabel metal2 33824 28616 33824 28616 0 gen_sym.Reg_Sym.data_out\[0\]
rlabel metal2 35896 30408 35896 30408 0 gen_sym.Reg_Sym.data_out\[1\]
rlabel metal2 33880 27384 33880 27384 0 mapper.bit_Q\[1\]
rlabel metal2 34720 29960 34720 29960 0 net1
rlabel metal2 55608 36120 55608 36120 0 net10
rlabel metal2 58184 48776 58184 48776 0 net100
rlabel metal2 55160 57610 55160 57610 0 net101
rlabel metal3 1246 41048 1246 41048 0 net102
rlabel metal3 58730 55832 58730 55832 0 net103
rlabel metal2 8232 55944 8232 55944 0 net104
rlabel metal2 58184 5544 58184 5544 0 net105
rlabel metal2 6776 2058 6776 2058 0 net106
rlabel metal2 58184 4984 58184 4984 0 net107
rlabel metal3 1246 30296 1246 30296 0 net108
rlabel metal2 49560 37968 49560 37968 0 net11
rlabel metal2 50456 40880 50456 40880 0 net12
rlabel metal2 51800 42448 51800 42448 0 net13
rlabel metal2 53032 44240 53032 44240 0 net14
rlabel metal2 53200 45752 53200 45752 0 net15
rlabel metal2 53928 51016 53928 51016 0 net16
rlabel metal2 53032 54432 53032 54432 0 net17
rlabel metal2 51576 54768 51576 54768 0 net18
rlabel metal2 40936 3976 40936 3976 0 net19
rlabel metal2 2072 26992 2072 26992 0 net2
rlabel metal2 55048 25928 55048 25928 0 net20
rlabel metal2 54264 27496 54264 27496 0 net21
rlabel metal3 48636 24136 48636 24136 0 net22
rlabel metal2 44184 4200 44184 4200 0 net23
rlabel metal2 48440 4200 48440 4200 0 net24
rlabel metal2 52080 6440 52080 6440 0 net25
rlabel metal2 54040 8680 54040 8680 0 net26
rlabel metal2 55944 12656 55944 12656 0 net27
rlabel metal2 54600 14448 54600 14448 0 net28
rlabel metal2 55272 17360 55272 17360 0 net29
rlabel metal2 27160 27944 27160 27944 0 net3
rlabel metal2 55160 20720 55160 20720 0 net30
rlabel metal2 54488 24248 54488 24248 0 net31
rlabel metal2 4312 29456 4312 29456 0 net32
rlabel metal2 4312 30688 4312 30688 0 net33
rlabel metal2 9128 31556 9128 31556 0 net34
rlabel metal2 4816 31528 4816 31528 0 net35
rlabel metal2 28504 29512 28504 29512 0 net36
rlabel metal2 30240 31192 30240 31192 0 net37
rlabel metal2 8008 23744 8008 23744 0 net38
rlabel metal2 9072 27608 9072 27608 0 net39
rlabel metal2 2072 25816 2072 25816 0 net4
rlabel metal3 8232 23688 8232 23688 0 net40
rlabel metal2 10136 23520 10136 23520 0 net41
rlabel metal2 15288 25816 15288 25816 0 net42
rlabel metal2 17864 24808 17864 24808 0 net43
rlabel metal2 33096 33768 33096 33768 0 net44
rlabel metal2 30072 28224 30072 28224 0 net45
rlabel metal3 33320 34104 33320 34104 0 net46
rlabel metal2 41720 31752 41720 31752 0 net47
rlabel metal2 38584 29008 38584 29008 0 net48
rlabel metal2 38024 27440 38024 27440 0 net49
rlabel metal2 9520 27832 9520 27832 0 net5
rlabel metal2 33376 27048 33376 27048 0 net50
rlabel metal2 17416 24024 17416 24024 0 net51
rlabel metal2 8792 23240 8792 23240 0 net52
rlabel metal2 30576 34888 30576 34888 0 net53
rlabel metal2 8904 32984 8904 32984 0 net54
rlabel metal2 8288 27944 8288 27944 0 net55
rlabel metal2 9576 30520 9576 30520 0 net56
rlabel metal2 9856 26936 9856 26936 0 net57
rlabel metal2 9688 27216 9688 27216 0 net58
rlabel metal2 28168 28112 28168 28112 0 net59
rlabel metal2 45416 35560 45416 35560 0 net6
rlabel metal2 38136 29680 38136 29680 0 net60
rlabel metal2 44520 28784 44520 28784 0 net61
rlabel metal2 44632 31920 44632 31920 0 net62
rlabel metal2 37240 27440 37240 27440 0 net63
rlabel metal2 28504 28224 28504 28224 0 net64
rlabel metal2 28392 29344 28392 29344 0 net65
rlabel metal2 12432 27160 12432 27160 0 net66
rlabel metal2 5992 29736 5992 29736 0 net67
rlabel metal2 11256 26488 11256 26488 0 net68
rlabel metal2 15008 26936 15008 26936 0 net69
rlabel metal2 48216 55776 48216 55776 0 net7
rlabel metal3 25816 28616 25816 28616 0 net70
rlabel metal3 1246 8792 1246 8792 0 net71
rlabel metal3 1246 53816 1246 53816 0 net72
rlabel metal2 58184 54768 58184 54768 0 net73
rlabel metal3 1246 28280 1246 28280 0 net74
rlabel metal3 58506 55160 58506 55160 0 net75
rlabel metal2 57736 3024 57736 3024 0 net76
rlabel metal2 58184 50960 58184 50960 0 net77
rlabel metal3 1470 29624 1470 29624 0 net78
rlabel metal3 53648 56280 53648 56280 0 net79
rlabel metal2 49448 53816 49448 53816 0 net8
rlabel metal3 58730 38360 58730 38360 0 net80
rlabel metal3 1246 37688 1246 37688 0 net81
rlabel metal2 5432 2030 5432 2030 0 net82
rlabel metal2 58240 39368 58240 39368 0 net83
rlabel metal2 58184 33040 58184 33040 0 net84
rlabel metal3 1246 18872 1246 18872 0 net85
rlabel metal2 58184 4256 58184 4256 0 net86
rlabel metal2 10248 56280 10248 56280 0 net87
rlabel metal2 58184 33936 58184 33936 0 net88
rlabel metal2 4760 2030 4760 2030 0 net89
rlabel metal2 48720 53368 48720 53368 0 net9
rlabel metal2 13608 56280 13608 56280 0 net90
rlabel metal2 58240 49896 58240 49896 0 net91
rlabel metal3 1246 16856 1246 16856 0 net92
rlabel metal3 58296 3304 58296 3304 0 net93
rlabel metal2 10920 56280 10920 56280 0 net94
rlabel metal2 54488 57778 54488 57778 0 net95
rlabel metal3 1246 32312 1246 32312 0 net96
rlabel metal2 58184 52752 58184 52752 0 net97
rlabel metal2 55048 56448 55048 56448 0 net98
rlabel metal2 7448 2030 7448 2030 0 net99
rlabel metal2 34832 36904 34832 36904 0 p_shaping_I.p_shaping_I.bit_in
rlabel metal2 38192 34328 38192 34328 0 p_shaping_I.p_shaping_I.bit_in_1
rlabel metal2 35112 34216 35112 34216 0 p_shaping_I.p_shaping_I.bit_in_2
rlabel metal2 44632 34048 44632 34048 0 p_shaping_I.p_shaping_I.counter\[0\]
rlabel metal2 37912 37296 37912 37296 0 p_shaping_I.p_shaping_I.counter\[1\]
rlabel metal2 40152 32368 40152 32368 0 p_shaping_I.p_shaping_I.ctl_1
rlabel metal2 36232 27832 36232 27832 0 p_shaping_Q.p_shaping_I.bit_in
rlabel metal2 38920 22568 38920 22568 0 p_shaping_Q.p_shaping_I.bit_in_1
rlabel metal2 42168 25368 42168 25368 0 p_shaping_Q.p_shaping_I.bit_in_2
rlabel metal2 43400 28840 43400 28840 0 p_shaping_Q.p_shaping_I.counter\[0\]
rlabel metal2 42168 22008 42168 22008 0 p_shaping_Q.p_shaping_I.counter\[1\]
rlabel metal2 40376 26600 40376 26600 0 p_shaping_Q.p_shaping_I.ctl_1
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
