VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OQPSK_RCOSINE_ALL
  CLASS BLOCK ;
  FOREIGN OQPSK_RCOSINE_ALL ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN ACK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 151.200 300.000 151.760 ;
    END
  END ACK
  PIN Bit_In
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END Bit_In
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END EN
  PIN I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 181.440 300.000 182.000 ;
    END
  END I[0]
  PIN I[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 296.000 239.120 300.000 ;
    END
  END I[10]
  PIN I[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 296.000 245.840 300.000 ;
    END
  END I[11]
  PIN I[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 296.000 242.480 300.000 ;
    END
  END I[12]
  PIN I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 178.080 300.000 178.640 ;
    END
  END I[1]
  PIN I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 188.160 300.000 188.720 ;
    END
  END I[2]
  PIN I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 201.600 300.000 202.160 ;
    END
  END I[3]
  PIN I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 208.320 300.000 208.880 ;
    END
  END I[4]
  PIN I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 218.400 300.000 218.960 ;
    END
  END I[5]
  PIN I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 235.200 300.000 235.760 ;
    END
  END I[6]
  PIN I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 255.360 300.000 255.920 ;
    END
  END I[7]
  PIN I[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 296.000 262.640 300.000 ;
    END
  END I[8]
  PIN I[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 296.000 255.920 300.000 ;
    END
  END I[9]
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 131.040 300.000 131.600 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 137.760 300.000 138.320 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 124.320 300.000 124.880 ;
    END
  END Q[12]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 0.000 242.480 4.000 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 43.680 300.000 44.240 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 60.480 300.000 61.040 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 73.920 300.000 74.480 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 87.360 300.000 87.920 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 104.160 300.000 104.720 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 120.960 300.000 121.520 ;
    END
  END Q[9]
  PIN REQ_SAMPLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END REQ_SAMPLE
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END RST
  PIN addI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END addI[0]
  PIN addI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END addI[1]
  PIN addI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END addI[2]
  PIN addI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END addI[3]
  PIN addI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END addI[4]
  PIN addI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 296.000 148.400 300.000 ;
    END
  END addI[5]
  PIN addQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END addQ[0]
  PIN addQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END addQ[1]
  PIN addQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END addQ[2]
  PIN addQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END addQ[3]
  PIN addQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END addQ[4]
  PIN addQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END addQ[5]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 241.920 300.000 242.480 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 272.160 300.000 272.720 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 275.520 300.000 276.080 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 13.440 300.000 14.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 248.640 300.000 249.200 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 296.000 266.000 300.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 191.520 300.000 192.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 296.000 276.080 300.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 194.880 300.000 195.440 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 164.640 300.000 165.200 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 20.160 300.000 20.720 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 296.000 50.960 300.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 168.000 300.000 168.560 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 296.000 67.760 300.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 245.280 300.000 245.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 16.800 300.000 17.360 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 296.000 54.320 300.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 296.000 272.720 300.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 262.080 300.000 262.640 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 296.000 269.360 300.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 278.880 300.000 279.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 296.000 40.880 300.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 26.880 300.000 27.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 23.520 300.000 24.080 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END io_oeb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 8.540 295.700 40.020 296.000 ;
        RECT 41.180 295.700 50.100 296.000 ;
        RECT 51.260 295.700 53.460 296.000 ;
        RECT 54.620 295.700 66.900 296.000 ;
        RECT 68.060 295.700 147.540 296.000 ;
        RECT 148.700 295.700 238.260 296.000 ;
        RECT 239.420 295.700 241.620 296.000 ;
        RECT 242.780 295.700 244.980 296.000 ;
        RECT 246.140 295.700 255.060 296.000 ;
        RECT 256.220 295.700 261.780 296.000 ;
        RECT 262.940 295.700 265.140 296.000 ;
        RECT 266.300 295.700 268.500 296.000 ;
        RECT 269.660 295.700 271.860 296.000 ;
        RECT 273.020 295.700 275.220 296.000 ;
        RECT 276.380 295.700 291.620 296.000 ;
        RECT 8.540 4.300 291.620 295.700 ;
        RECT 8.540 4.000 23.220 4.300 ;
        RECT 24.380 4.000 26.580 4.300 ;
        RECT 27.740 4.000 33.300 4.300 ;
        RECT 34.460 4.000 36.660 4.300 ;
        RECT 37.820 4.000 204.660 4.300 ;
        RECT 205.820 4.000 218.100 4.300 ;
        RECT 219.260 4.000 241.620 4.300 ;
        RECT 242.780 4.000 258.420 4.300 ;
        RECT 259.580 4.000 291.620 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 279.740 296.660 286.020 ;
        RECT 4.000 278.580 295.700 279.740 ;
        RECT 4.000 276.380 296.660 278.580 ;
        RECT 4.000 275.220 295.700 276.380 ;
        RECT 4.000 273.020 296.660 275.220 ;
        RECT 4.000 271.860 295.700 273.020 ;
        RECT 4.000 269.660 296.660 271.860 ;
        RECT 4.300 268.500 296.660 269.660 ;
        RECT 4.000 262.940 296.660 268.500 ;
        RECT 4.000 261.780 295.700 262.940 ;
        RECT 4.000 256.220 296.660 261.780 ;
        RECT 4.000 255.060 295.700 256.220 ;
        RECT 4.000 249.500 296.660 255.060 ;
        RECT 4.000 248.340 295.700 249.500 ;
        RECT 4.000 246.140 296.660 248.340 ;
        RECT 4.000 244.980 295.700 246.140 ;
        RECT 4.000 242.780 296.660 244.980 ;
        RECT 4.000 241.620 295.700 242.780 ;
        RECT 4.000 236.060 296.660 241.620 ;
        RECT 4.000 234.900 295.700 236.060 ;
        RECT 4.000 219.260 296.660 234.900 ;
        RECT 4.000 218.100 295.700 219.260 ;
        RECT 4.000 209.180 296.660 218.100 ;
        RECT 4.000 208.020 295.700 209.180 ;
        RECT 4.000 205.820 296.660 208.020 ;
        RECT 4.300 204.660 296.660 205.820 ;
        RECT 4.000 202.460 296.660 204.660 ;
        RECT 4.000 201.300 295.700 202.460 ;
        RECT 4.000 195.740 296.660 201.300 ;
        RECT 4.000 194.580 295.700 195.740 ;
        RECT 4.000 192.380 296.660 194.580 ;
        RECT 4.000 191.220 295.700 192.380 ;
        RECT 4.000 189.020 296.660 191.220 ;
        RECT 4.300 187.860 295.700 189.020 ;
        RECT 4.000 182.300 296.660 187.860 ;
        RECT 4.000 181.140 295.700 182.300 ;
        RECT 4.000 178.940 296.660 181.140 ;
        RECT 4.000 177.780 295.700 178.940 ;
        RECT 4.000 168.860 296.660 177.780 ;
        RECT 4.300 167.700 295.700 168.860 ;
        RECT 4.000 165.500 296.660 167.700 ;
        RECT 4.300 164.340 295.700 165.500 ;
        RECT 4.000 162.140 296.660 164.340 ;
        RECT 4.300 160.980 296.660 162.140 ;
        RECT 4.000 158.780 296.660 160.980 ;
        RECT 4.300 157.620 296.660 158.780 ;
        RECT 4.000 155.420 296.660 157.620 ;
        RECT 4.300 154.260 296.660 155.420 ;
        RECT 4.000 152.060 296.660 154.260 ;
        RECT 4.300 150.900 295.700 152.060 ;
        RECT 4.000 148.700 296.660 150.900 ;
        RECT 4.300 147.540 296.660 148.700 ;
        RECT 4.000 145.340 296.660 147.540 ;
        RECT 4.300 144.180 296.660 145.340 ;
        RECT 4.000 141.980 296.660 144.180 ;
        RECT 4.300 140.820 296.660 141.980 ;
        RECT 4.000 138.620 296.660 140.820 ;
        RECT 4.300 137.460 295.700 138.620 ;
        RECT 4.000 135.260 296.660 137.460 ;
        RECT 4.300 134.100 296.660 135.260 ;
        RECT 4.000 131.900 296.660 134.100 ;
        RECT 4.300 130.740 295.700 131.900 ;
        RECT 4.000 128.540 296.660 130.740 ;
        RECT 4.300 127.380 296.660 128.540 ;
        RECT 4.000 125.180 296.660 127.380 ;
        RECT 4.300 124.020 295.700 125.180 ;
        RECT 4.000 121.820 296.660 124.020 ;
        RECT 4.300 120.660 295.700 121.820 ;
        RECT 4.000 118.460 296.660 120.660 ;
        RECT 4.300 117.300 296.660 118.460 ;
        RECT 4.000 115.100 296.660 117.300 ;
        RECT 4.300 113.940 296.660 115.100 ;
        RECT 4.000 111.740 296.660 113.940 ;
        RECT 4.300 110.580 296.660 111.740 ;
        RECT 4.000 108.380 296.660 110.580 ;
        RECT 4.300 107.220 296.660 108.380 ;
        RECT 4.000 105.020 296.660 107.220 ;
        RECT 4.000 103.860 295.700 105.020 ;
        RECT 4.000 94.940 296.660 103.860 ;
        RECT 4.300 93.780 296.660 94.940 ;
        RECT 4.000 88.220 296.660 93.780 ;
        RECT 4.000 87.060 295.700 88.220 ;
        RECT 4.000 84.860 296.660 87.060 ;
        RECT 4.300 83.700 296.660 84.860 ;
        RECT 4.000 74.780 296.660 83.700 ;
        RECT 4.000 73.620 295.700 74.780 ;
        RECT 4.000 61.340 296.660 73.620 ;
        RECT 4.000 60.180 295.700 61.340 ;
        RECT 4.000 44.540 296.660 60.180 ;
        RECT 4.300 43.380 295.700 44.540 ;
        RECT 4.000 27.740 296.660 43.380 ;
        RECT 4.000 26.580 295.700 27.740 ;
        RECT 4.000 24.380 296.660 26.580 ;
        RECT 4.000 23.220 295.700 24.380 ;
        RECT 4.000 21.020 296.660 23.220 ;
        RECT 4.000 19.860 295.700 21.020 ;
        RECT 4.000 17.660 296.660 19.860 ;
        RECT 4.000 16.500 295.700 17.660 ;
        RECT 4.000 14.300 296.660 16.500 ;
        RECT 4.000 13.140 295.700 14.300 ;
        RECT 4.000 6.860 296.660 13.140 ;
      LAYER Metal4 ;
        RECT 39.900 282.840 232.820 286.070 ;
        RECT 39.900 15.080 98.740 282.840 ;
        RECT 100.940 15.080 175.540 282.840 ;
        RECT 177.740 15.080 232.820 282.840 ;
        RECT 39.900 6.810 232.820 15.080 ;
  END
END OQPSK_RCOSINE_ALL
END LIBRARY

