// This is the unpowered netlist.
module OQPSK_RCOSINE_ALL (ACK,
    Bit_In,
    EN,
    REQ_SAMPLE,
    RST,
    I,
    Q,
    addI,
    addQ,
    io_oeb);
 input ACK;
 input Bit_In;
 input EN;
 input REQ_SAMPLE;
 input RST;
 output [12:0] I;
 output [12:0] Q;
 output [5:0] addI;
 output [5:0] addQ;
 output [37:0] io_oeb;

 wire net100;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net101;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net102;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net71;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire \gen_sym.Reg_2M.data_in ;
 wire \gen_sym.Reg_2M.data_out ;
 wire \gen_sym.Reg_2M.enable ;
 wire \gen_sym.Reg_Sym.data_out[0] ;
 wire \gen_sym.Reg_Sym.data_out[1] ;
 wire \mapper.bit_Q[1] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net8;
 wire net9;
 wire \p_shaping_I.p_shaping_I.bit_in ;
 wire \p_shaping_I.p_shaping_I.bit_in_1 ;
 wire \p_shaping_I.p_shaping_I.bit_in_2 ;
 wire \p_shaping_I.p_shaping_I.counter[0] ;
 wire \p_shaping_I.p_shaping_I.counter[1] ;
 wire \p_shaping_I.p_shaping_I.ctl_1 ;
 wire \p_shaping_Q.p_shaping_I.bit_in ;
 wire \p_shaping_Q.p_shaping_I.bit_in_1 ;
 wire \p_shaping_Q.p_shaping_I.bit_in_2 ;
 wire \p_shaping_Q.p_shaping_I.counter[0] ;
 wire \p_shaping_Q.p_shaping_I.counter[1] ;
 wire \p_shaping_Q.p_shaping_I.ctl_1 ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1381__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A2 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A1 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__B1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A4 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1436__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__I (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__B (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__B2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__C (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A3 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__I (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__I (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A3 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__B (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A3 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1572__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__B1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__C (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I0 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__I (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__I (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__B2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__B (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__I0 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__B (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__B (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__B (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__B (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__B (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A3 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A3 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__B1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__B2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A3 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__B (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__B (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__B (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__B (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__B (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__B (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__B (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__B2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__B (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__B (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__B (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__B1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__C (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__B (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__B (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__I (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__B (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__B (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__B (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A3 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__B (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__B (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__B (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A3 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A3 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__B2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__B (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A3 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__C (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__B (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__B2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__B (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A3 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__B2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A3 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A4 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__B2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__C2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__S0 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A3 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A4 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A3 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__B2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__B2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__B (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__B (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__B2 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__C (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__B (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__C (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__B2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__B2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__S (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__B (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__B (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__C (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__C (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__B1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__B2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__I (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__C (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__B (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__B (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A3 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__C (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__B2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__B1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__B (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A3 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__I (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__B (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__B (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__B (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__B (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__B (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A3 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A1 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__B (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A3 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A2 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__B2 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__C (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__B1 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__C1 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A3 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__B (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__B (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__C (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__B1 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A3 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A3 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A4 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__B1 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A3 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__S (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A3 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__I0 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A4 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__B (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__B (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__B (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__I (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A3 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__B1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__B (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__C (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A3 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__C (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A3 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__I (.I(\p_shaping_I.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A3 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A4 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__B (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__B1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__C (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__B2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A1 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__D (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__D (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(\p_shaping_I.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ACK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(Bit_In));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(EN));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(REQ_SAMPLE));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(RST));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_100 (.Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_101 (.Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_102 (.Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_103 (.Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_104 (.Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_105 (.Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_106 (.Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_107 (.Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__tieh OQPSK_RCOSINE_ALL_108 (.Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel OQPSK_RCOSINE_ALL_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1373_ (.I(net35),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1374_ (.I(_1200_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1375_ (.I(_1211_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1376_ (.I(_1220_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1377_ (.I(net54),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1378_ (.I(_1241_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1379_ (.I(_1252_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1380_ (.I(_1263_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1381_ (.I(net35),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1382_ (.I(_1285_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1383_ (.I(net54),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1384_ (.I(_1307_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1385_ (.A1(_1296_),
    .A2(_1318_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1386_ (.I(_1200_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1387_ (.I(net33),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1388_ (.I(_1350_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1389_ (.I(net32),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1390_ (.I(_1372_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1391_ (.A1(_1361_),
    .A2(_0032_),
    .A3(_1307_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1392_ (.A1(_1339_),
    .A2(_0043_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1393_ (.I(net36),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1394_ (.I(_0065_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1395_ (.I(net53),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1396_ (.A1(_0076_),
    .A2(_0087_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1397_ (.A1(_1328_),
    .A2(_0054_),
    .B(_0098_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1398_ (.I(net53),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1399_ (.I(net33),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1400_ (.I(net54),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1401_ (.A1(_0129_),
    .A2(_0140_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1402_ (.I(_0151_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1403_ (.I(net36),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1404_ (.A1(_1296_),
    .A2(_0162_),
    .B(_0173_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1405_ (.A1(_1296_),
    .A2(_0151_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1406_ (.I(_0065_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1407_ (.I(net53),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1408_ (.A1(_0205_),
    .A2(_0216_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1409_ (.A1(_0118_),
    .A2(_0183_),
    .B1(_0194_),
    .B2(_0227_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1410_ (.A1(_0107_),
    .A2(_0237_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1411_ (.I(_1361_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1412_ (.I(_1372_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1413_ (.I(_0270_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1414_ (.I(_0281_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1415_ (.A1(_0259_),
    .A2(_0291_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1416_ (.A1(_1230_),
    .A2(_1274_),
    .A3(_0248_),
    .A4(_0302_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1417_ (.I(_0313_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1418_ (.I(_0324_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1419_ (.I(net39),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1420_ (.I(_0344_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1421_ (.I(_0355_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1422_ (.I(net38),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1423_ (.I(_0377_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1424_ (.I(_0387_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1425_ (.I(net41),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1426_ (.I(_0409_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1427_ (.I(net52),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1428_ (.I(_0430_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1429_ (.A1(_0366_),
    .A2(_0398_),
    .A3(_0419_),
    .A4(_0441_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1430_ (.I(_0409_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1431_ (.I(net39),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1432_ (.I(_0472_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1433_ (.I(net52),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1434_ (.A1(_0483_),
    .A2(_0387_),
    .A3(_0493_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1435_ (.I(net41),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1436_ (.A1(_0508_),
    .A2(_0493_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1437_ (.I(net42),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1438_ (.A1(_0462_),
    .A2(_0500_),
    .B(_0515_),
    .C(_0524_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1439_ (.I(net42),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1440_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1441_ (.A1(_0483_),
    .A2(_0508_),
    .A3(_0493_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1442_ (.A1(_0530_),
    .A2(_0531_),
    .B(net51),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1443_ (.I(_0472_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1444_ (.I(net52),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1445_ (.I(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1446_ (.I(net41),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1447_ (.A1(_0533_),
    .A2(_0535_),
    .B(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1448_ (.I(net51),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1449_ (.A1(_0530_),
    .A2(_0537_),
    .B(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1450_ (.A1(_0528_),
    .A2(_0532_),
    .B(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1451_ (.A1(_0451_),
    .A2(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1452_ (.I(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1453_ (.I(_0542_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1454_ (.I(net1),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1455_ (.A1(\gen_sym.Reg_Sym.data_out[1] ),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1456_ (.I(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1457_ (.I(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1458_ (.I(_0546_),
    .Z(\p_shaping_I.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1459_ (.A1(_0543_),
    .A2(\gen_sym.Reg_Sym.data_out[0] ),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1460_ (.I(_0547_),
    .Z(\mapper.bit_Q[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1461_ (.I(net44),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1462_ (.I(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1463_ (.I(_0313_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1464_ (.I(net60),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1465_ (.I(_0544_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1466_ (.A1(\p_shaping_I.p_shaping_I.ctl_1 ),
    .A2(_0551_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1467_ (.A1(_0551_),
    .A2(_0552_),
    .B(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1468_ (.A1(_0550_),
    .A2(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1469_ (.A1(_0549_),
    .A2(_0550_),
    .B(_0555_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1470_ (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1471_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1472_ (.I(\p_shaping_Q.p_shaping_I.bit_in ),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1473_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1474_ (.A1(net61),
    .A2(\p_shaping_Q.p_shaping_I.ctl_1 ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1475_ (.A1(_0551_),
    .A2(_0559_),
    .B(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1476_ (.A1(_0542_),
    .A2(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1477_ (.A1(_0557_),
    .A2(net48),
    .B(_0562_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1478_ (.A1(net3),
    .A2(net2),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1479_ (.I(_0563_),
    .Z(\gen_sym.Reg_2M.data_in ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1480_ (.A1(net45),
    .A2(_0542_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1481_ (.I(_0564_),
    .Z(\gen_sym.Reg_2M.enable ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1482_ (.I(_0551_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1483_ (.A1(_0565_),
    .A2(net46),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1484_ (.A1(_0565_),
    .A2(net48),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1485_ (.I(\p_shaping_Q.p_shaping_I.counter[1] ),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1486_ (.I(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1487_ (.I(_0508_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1488_ (.I(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1489_ (.I(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1490_ (.I(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1491_ (.I(net38),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1492_ (.A1(_0344_),
    .A2(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1493_ (.I(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1494_ (.I(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1495_ (.I(_0534_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1496_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1497_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1498_ (.I(_0568_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1499_ (.I(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1500_ (.I(net51),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1501_ (.I(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1502_ (.A1(_0580_),
    .A2(_0582_),
    .B(_0575_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1503_ (.I(_0377_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1504_ (.I(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1505_ (.I(_0493_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1506_ (.A1(_0585_),
    .A2(_0586_),
    .B(_0462_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1507_ (.I(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1508_ (.I(_0483_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1509_ (.I(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1510_ (.I(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1511_ (.I(_0524_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1512_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1513_ (.A1(_0578_),
    .A2(_0583_),
    .B1(_0588_),
    .B2(_0591_),
    .C(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1514_ (.I(_0377_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1515_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1516_ (.I(_0534_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1517_ (.A1(_0533_),
    .A2(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1518_ (.I(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1519_ (.A1(_0596_),
    .A2(_0579_),
    .A3(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1520_ (.I(_0409_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1521_ (.I(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1522_ (.I(_0441_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1523_ (.A1(_0344_),
    .A2(_0572_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1524_ (.I(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1525_ (.I(_0605_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1526_ (.A1(_0602_),
    .A2(_0603_),
    .A3(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1527_ (.A1(_0593_),
    .A2(_0600_),
    .A3(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1528_ (.I(_0536_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1529_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1530_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1531_ (.I(_0524_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1532_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1533_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1534_ (.I(net43),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1535_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1536_ (.A1(_0611_),
    .A2(_0614_),
    .B(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1537_ (.A1(_0571_),
    .A2(_0575_),
    .B1(_0594_),
    .B2(_0608_),
    .C(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1538_ (.A1(_0567_),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1539_ (.I(_0538_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1540_ (.A1(_0533_),
    .A2(_0387_),
    .A3(_0536_),
    .A4(_0597_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1541_ (.A1(_0612_),
    .A2(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1542_ (.A1(_0620_),
    .A2(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1543_ (.I(_0344_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1544_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1545_ (.I(_0430_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1546_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1547_ (.A1(_0625_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1548_ (.I(_0355_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1549_ (.I(_0535_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1550_ (.I(_0462_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1551_ (.A1(_0629_),
    .A2(_0630_),
    .B(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1552_ (.I(_0624_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1553_ (.I(_0626_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1554_ (.A1(_0633_),
    .A2(_0569_),
    .A3(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1555_ (.A1(_0628_),
    .A2(_0632_),
    .B(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1556_ (.A1(_0483_),
    .A2(_0572_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1557_ (.A1(_0627_),
    .A2(_0637_),
    .B(_0631_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1558_ (.I(_0584_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1559_ (.A1(_0633_),
    .A2(_0639_),
    .B(_0630_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1560_ (.I(_0529_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1561_ (.I(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1562_ (.A1(net39),
    .A2(net38),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1563_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1564_ (.A1(_0579_),
    .A2(_0599_),
    .A3(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1565_ (.A1(_0638_),
    .A2(_0640_),
    .B(_0642_),
    .C(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1566_ (.A1(_0601_),
    .A2(_0598_),
    .A3(_0574_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1567_ (.I(_0572_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1568_ (.A1(_0648_),
    .A2(_0536_),
    .A3(_0535_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1569_ (.A1(_0612_),
    .A2(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1570_ (.I(_0581_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1571_ (.A1(_0647_),
    .A2(_0650_),
    .B(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1572_ (.A1(_0623_),
    .A2(_0636_),
    .B1(_0646_),
    .B2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1573_ (.A1(\p_shaping_Q.p_shaping_I.counter[0] ),
    .A2(\p_shaping_Q.p_shaping_I.counter[1] ),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1574_ (.I(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1575_ (.I(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1576_ (.A1(_0653_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1577_ (.I(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1578_ (.I(_0419_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1579_ (.A1(_0648_),
    .A2(_0576_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1580_ (.A1(_0630_),
    .A2(_0644_),
    .B(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1581_ (.A1(_0629_),
    .A2(_0596_),
    .B(_0660_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1582_ (.A1(_0659_),
    .A2(_0661_),
    .A3(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1583_ (.I(_0508_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _1584_ (.I0(_0387_),
    .I1(_0533_),
    .S(_0534_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1585_ (.A1(_0664_),
    .A2(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1586_ (.I(_0597_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1587_ (.A1(_0398_),
    .A2(_0667_),
    .B(_0664_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1588_ (.I(_0530_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1589_ (.A1(_0605_),
    .A2(_0666_),
    .B1(_0668_),
    .B2(_0669_),
    .C(_0615_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1590_ (.I0(_0605_),
    .I1(_0644_),
    .S(_0626_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1591_ (.I(_0597_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1592_ (.A1(_0366_),
    .A2(_0601_),
    .A3(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1593_ (.A1(_0659_),
    .A2(_0671_),
    .B(_0673_),
    .C(_0669_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1594_ (.I(_0620_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1595_ (.I(_0524_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1596_ (.A1(_0676_),
    .A2(_0531_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1597_ (.A1(_0675_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1598_ (.A1(_0663_),
    .A2(_0670_),
    .B1(_0674_),
    .B2(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1599_ (.I(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1600_ (.A1(_0658_),
    .A2(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1601_ (.A1(_0619_),
    .A2(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1602_ (.I(_0682_),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1603_ (.A1(_0658_),
    .A2(_0680_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1604_ (.A1(_0619_),
    .A2(_0681_),
    .B(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1605_ (.I(_0584_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1606_ (.I(_0462_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1607_ (.A1(_0633_),
    .A2(_0685_),
    .B(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1608_ (.A1(_0628_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1609_ (.I(_0676_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(_0689_),
    .A2(_0537_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1611_ (.A1(_0590_),
    .A2(_0685_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1612_ (.I(_0500_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1613_ (.A1(_0579_),
    .A2(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1614_ (.A1(_0602_),
    .A2(_0691_),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1615_ (.A1(_0530_),
    .A2(_0538_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1616_ (.I(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1617_ (.I(_0568_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1618_ (.A1(_0589_),
    .A2(_0672_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1619_ (.A1(_0472_),
    .A2(_0377_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1620_ (.I(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1621_ (.A1(_0697_),
    .A2(_0698_),
    .A3(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1622_ (.A1(_0613_),
    .A2(_0666_),
    .A3(_0701_),
    .B(_0651_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1623_ (.A1(_0688_),
    .A2(_0690_),
    .B1(_0694_),
    .B2(_0696_),
    .C(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1624_ (.I(\p_shaping_Q.p_shaping_I.bit_in ),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1625_ (.A1(_0704_),
    .A2(_0680_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1626_ (.A1(_0703_),
    .A2(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1627_ (.I(_0654_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1628_ (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1629_ (.A1(_0603_),
    .A2(_0574_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1630_ (.A1(_0366_),
    .A2(_0398_),
    .B(_0586_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1631_ (.A1(_0709_),
    .A2(_0710_),
    .B(_0610_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1632_ (.A1(_0596_),
    .A2(_0627_),
    .B(_0569_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1633_ (.A1(_0592_),
    .A2(_0615_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1634_ (.A1(_0712_),
    .A2(_0640_),
    .B(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1635_ (.A1(_0625_),
    .A2(_0441_),
    .B(_0609_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1636_ (.A1(_0641_),
    .A2(_0581_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1637_ (.A1(_0715_),
    .A2(_0693_),
    .B(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1638_ (.A1(_0624_),
    .A2(_0595_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1639_ (.I0(_0718_),
    .I1(_0699_),
    .S(_0626_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1640_ (.I(_0568_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1641_ (.A1(_0720_),
    .A2(_0599_),
    .B(_0669_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1642_ (.A1(_0642_),
    .A2(_0531_),
    .B1(_0719_),
    .B2(_0721_),
    .C(_0651_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1643_ (.A1(_0711_),
    .A2(_0714_),
    .B(_0717_),
    .C(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1644_ (.A1(_0708_),
    .A2(_0653_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1645_ (.I(_0643_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1646_ (.A1(_0472_),
    .A2(net40),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1647_ (.I(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1648_ (.A1(_0419_),
    .A2(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1649_ (.A1(_0586_),
    .A2(_0604_),
    .B(_0664_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1650_ (.A1(_0355_),
    .A2(_0595_),
    .B(_0430_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1651_ (.A1(_0725_),
    .A2(_0728_),
    .B1(_0729_),
    .B2(_0730_),
    .C(_0592_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1652_ (.A1(_0647_),
    .A2(_0650_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1653_ (.A1(_0592_),
    .A2(_0621_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1654_ (.A1(_0651_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1655_ (.I(_0576_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1656_ (.A1(_0629_),
    .A2(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1657_ (.A1(_0366_),
    .A2(_0601_),
    .A3(_0630_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1658_ (.A1(_0736_),
    .A2(_0715_),
    .B(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _1659_ (.A1(_0582_),
    .A2(_0731_),
    .A3(_0732_),
    .B1(_0734_),
    .B2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1660_ (.A1(_0672_),
    .A2(_0718_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1661_ (.A1(_0589_),
    .A2(_0585_),
    .B(_0441_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1662_ (.A1(_0740_),
    .A2(_0741_),
    .B(_0659_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1663_ (.I(_0730_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1664_ (.A1(_0587_),
    .A2(_0743_),
    .B(_0695_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1665_ (.A1(_0720_),
    .A2(_0692_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1666_ (.A1(_0676_),
    .A2(_0620_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1667_ (.A1(_0632_),
    .A2(_0745_),
    .B(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1668_ (.A1(_0624_),
    .A2(_0648_),
    .B(_0576_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1669_ (.A1(_0735_),
    .A2(_0699_),
    .B(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1670_ (.A1(_0631_),
    .A2(_0727_),
    .B(_0676_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1671_ (.A1(_0749_),
    .A2(_0750_),
    .B(_0532_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1672_ (.A1(_0742_),
    .A2(_0744_),
    .B(_0747_),
    .C(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1673_ (.A1(_0556_),
    .A2(_0739_),
    .A3(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1674_ (.A1(_0707_),
    .A2(_0724_),
    .A3(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1675_ (.A1(_0706_),
    .A2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1676_ (.I(\p_shaping_Q.p_shaping_I.counter[1] ),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1677_ (.I(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1678_ (.A1(_0757_),
    .A2(_0618_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1679_ (.A1(_0625_),
    .A2(_0639_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1680_ (.I(_0355_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1681_ (.I(_0735_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1682_ (.A1(_0760_),
    .A2(_0580_),
    .A3(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1683_ (.I(_0648_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1684_ (.A1(_0611_),
    .A2(_0578_),
    .A3(_0759_),
    .B1(_0762_),
    .B2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1685_ (.I(_0686_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1686_ (.A1(_0419_),
    .A2(_0667_),
    .A3(_0605_),
    .A4(_0573_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1687_ (.I(_0642_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1688_ (.A1(_0765_),
    .A2(_0665_),
    .B(_0766_),
    .C(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1689_ (.I(_0580_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1690_ (.I(_0725_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1691_ (.A1(_0767_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1692_ (.I(_0582_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1693_ (.A1(_0769_),
    .A2(_0771_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1694_ (.A1(_0623_),
    .A2(_0764_),
    .B1(_0768_),
    .B2(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1695_ (.A1(_0758_),
    .A2(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1696_ (.A1(_0756_),
    .A2(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1697_ (.A1(_0755_),
    .A2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1698_ (.A1(_0684_),
    .A2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1699_ (.A1(_0724_),
    .A2(_0753_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1700_ (.A1(_0656_),
    .A2(_0706_),
    .A3(_0779_),
    .B1(_0755_),
    .B2(_0776_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1701_ (.I(_0637_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1702_ (.A1(_0634_),
    .A2(_0781_),
    .B(_0697_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1703_ (.A1(_0634_),
    .A2(_0644_),
    .B(_0615_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1704_ (.I(_0641_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1705_ (.A1(_0782_),
    .A2(_0783_),
    .B(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1706_ (.A1(_0760_),
    .A2(_0763_),
    .A3(_0686_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1707_ (.A1(_0569_),
    .A2(_0781_),
    .B1(_0727_),
    .B2(_0639_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1708_ (.A1(_0786_),
    .A2(_0787_),
    .B(_0675_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1709_ (.A1(_0409_),
    .A2(_0726_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1710_ (.A1(_0685_),
    .A2(_0698_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1711_ (.A1(_0789_),
    .A2(_0790_),
    .B(_0695_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1712_ (.A1(_0785_),
    .A2(_0788_),
    .A3(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1713_ (.A1(_0680_),
    .A2(_0703_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1714_ (.A1(_0704_),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1715_ (.A1(_0792_),
    .A2(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1716_ (.A1(_0558_),
    .A2(_0560_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1717_ (.A1(_0541_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1718_ (.A1(_0625_),
    .A2(_0639_),
    .A3(_0609_),
    .A4(_0672_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1719_ (.A1(_0669_),
    .A2(_0798_),
    .B(_0766_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1720_ (.A1(_0595_),
    .A2(_0535_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1721_ (.A1(_0641_),
    .A2(_0581_),
    .B(_0800_),
    .C(_0664_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1722_ (.A1(_0585_),
    .A2(_0612_),
    .A3(_0620_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1723_ (.A1(_0633_),
    .A2(_0801_),
    .B1(_0802_),
    .B2(_0789_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1724_ (.A1(_0586_),
    .A2(_0699_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1725_ (.A1(_0800_),
    .A2(_0804_),
    .B(_0695_),
    .C(_0720_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1726_ (.A1(_0582_),
    .A2(_0799_),
    .B(_0803_),
    .C(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1727_ (.A1(_0653_),
    .A2(_0723_),
    .B(_0708_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1728_ (.A1(_0797_),
    .A2(_0806_),
    .A3(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1729_ (.A1(_0655_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1730_ (.A1(_0618_),
    .A2(_0774_),
    .B(_0757_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1731_ (.A1(_0689_),
    .A2(_0675_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1732_ (.I(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1733_ (.A1(_0611_),
    .A2(_0743_),
    .B(_0649_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1734_ (.I(_0660_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1735_ (.I(_0602_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1736_ (.A1(_0759_),
    .A2(_0515_),
    .B1(_0814_),
    .B2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1737_ (.I(_0627_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1738_ (.I(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1739_ (.I(_0760_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1740_ (.A1(_0819_),
    .A2(_0763_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1741_ (.A1(_0818_),
    .A2(_0820_),
    .B(_0696_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1742_ (.I(_0781_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1743_ (.I(_0609_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1744_ (.A1(_0823_),
    .A2(_0817_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1745_ (.I(_0667_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1746_ (.A1(_0825_),
    .A2(_0822_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1747_ (.A1(_0822_),
    .A2(_0824_),
    .B1(_0826_),
    .B2(_0687_),
    .C(_0746_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1748_ (.A1(_0812_),
    .A2(_0813_),
    .B1(_0816_),
    .B2(_0821_),
    .C(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1749_ (.A1(_0810_),
    .A2(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1750_ (.A1(_0566_),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1751_ (.A1(_0795_),
    .A2(_0809_),
    .A3(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1752_ (.A1(_0778_),
    .A2(_0780_),
    .A3(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1753_ (.I(_0832_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1754_ (.A1(_0780_),
    .A2(_0831_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1755_ (.A1(_0780_),
    .A2(_0831_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1756_ (.A1(_0684_),
    .A2(_0777_),
    .A3(_0833_),
    .B(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1757_ (.A1(_0795_),
    .A2(_0809_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1758_ (.A1(_0656_),
    .A2(_0795_),
    .A3(_0808_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1759_ (.A1(_0836_),
    .A2(_0830_),
    .B(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1760_ (.I(_0570_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1761_ (.A1(_0578_),
    .A2(_0770_),
    .B(_0692_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1762_ (.A1(_0666_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1763_ (.I(_0784_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1764_ (.A1(_0839_),
    .A2(_0665_),
    .B(_0841_),
    .C(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1765_ (.A1(_0629_),
    .A2(_0577_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1766_ (.A1(_0571_),
    .A2(_0844_),
    .A3(_0741_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1767_ (.A1(_0591_),
    .A2(_0817_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1768_ (.I(_0710_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1769_ (.A1(_0765_),
    .A2(_0575_),
    .B1(_0846_),
    .B2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1770_ (.I(_0593_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1771_ (.A1(_0845_),
    .A2(_0848_),
    .B(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1772_ (.I(_0772_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1773_ (.A1(_0843_),
    .A2(_0850_),
    .B(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1774_ (.I(_0761_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1775_ (.A1(_0763_),
    .A2(_0761_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1776_ (.A1(_0853_),
    .A2(_0770_),
    .B(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1777_ (.A1(_0688_),
    .A2(_0855_),
    .B(_0812_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1778_ (.A1(_0688_),
    .A2(_0855_),
    .B(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1779_ (.A1(_0852_),
    .A2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1780_ (.I(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1781_ (.A1(_0618_),
    .A2(_0774_),
    .A3(_0828_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1782_ (.A1(_0859_),
    .A2(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1783_ (.A1(_0858_),
    .A2(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1784_ (.A1(_0567_),
    .A2(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1785_ (.I(_0704_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1786_ (.A1(_0792_),
    .A2(_0793_),
    .B(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1787_ (.I(_0686_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1788_ (.A1(_0577_),
    .A2(_0700_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1789_ (.A1(_0725_),
    .A2(_0668_),
    .B(_0642_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1790_ (.A1(_0866_),
    .A2(_0867_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1791_ (.I(_0451_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1792_ (.A1(_0616_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1793_ (.A1(_0823_),
    .A2(_0847_),
    .B(_0713_),
    .C(_0600_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1794_ (.A1(_0610_),
    .A2(_0574_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1795_ (.A1(_0589_),
    .A2(_0398_),
    .A3(_0667_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1796_ (.A1(_0588_),
    .A2(_0873_),
    .B(_0874_),
    .C(_0716_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1797_ (.A1(_0869_),
    .A2(_0871_),
    .B(_0872_),
    .C(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1798_ (.A1(_0865_),
    .A2(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1799_ (.A1(_0739_),
    .A2(_0752_),
    .A3(_0806_),
    .B(_0556_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1800_ (.A1(_0825_),
    .A2(_0700_),
    .B(_0748_),
    .C(_0610_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1801_ (.A1(_0733_),
    .A2(_0673_),
    .A3(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1802_ (.A1(_0616_),
    .A2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1803_ (.A1(_0760_),
    .A2(_0634_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1804_ (.A1(_0882_),
    .A2(_0804_),
    .B(_0602_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1805_ (.A1(_0823_),
    .A2(_0844_),
    .A3(_0741_),
    .B(_0784_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1806_ (.I(_0675_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1807_ (.A1(_0823_),
    .A2(_0814_),
    .B(_0600_),
    .C(_0689_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1808_ (.A1(_0883_),
    .A2(_0884_),
    .B(_0885_),
    .C(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1809_ (.A1(_0881_),
    .A2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1810_ (.A1(_0878_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1811_ (.I(_0707_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1812_ (.A1(_0797_),
    .A2(_0889_),
    .B(_0007_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1813_ (.A1(_0541_),
    .A2(_0796_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1814_ (.I(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1815_ (.I(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1816_ (.A1(_0878_),
    .A2(_0888_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1817_ (.A1(_0893_),
    .A2(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1818_ (.A1(_0877_),
    .A2(_0890_),
    .A3(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1819_ (.I(_0890_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1820_ (.A1(_0897_),
    .A2(_0895_),
    .B(_0877_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1821_ (.A1(_0896_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1822_ (.A1(_0838_),
    .A2(_0863_),
    .A3(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1823_ (.A1(_0835_),
    .A2(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1824_ (.I(_0901_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1825_ (.A1(_0852_),
    .A2(_0857_),
    .A3(_0860_),
    .B(_0859_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1826_ (.I(_0616_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1827_ (.A1(_0817_),
    .A2(_0770_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1828_ (.A1(_0854_),
    .A2(_0904_),
    .B(_0815_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1829_ (.I(_0585_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1830_ (.I(_0727_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1831_ (.A1(_0906_),
    .A2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1832_ (.A1(_0537_),
    .A2(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1833_ (.A1(_0614_),
    .A2(_0905_),
    .A3(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1834_ (.A1(_0839_),
    .A2(_0822_),
    .B(_0721_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1835_ (.I(_0767_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1836_ (.I(_0606_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1837_ (.A1(_0853_),
    .A2(_0913_),
    .B(_0575_),
    .C(_0769_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1838_ (.A1(_0912_),
    .A2(_0903_),
    .A3(_0766_),
    .A4(_0914_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _1839_ (.A1(_0903_),
    .A2(_0910_),
    .A3(_0911_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1840_ (.A1(_0902_),
    .A2(_0916_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1841_ (.A1(_0567_),
    .A2(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1842_ (.A1(_0679_),
    .A2(_0703_),
    .A3(_0792_),
    .A4(_0876_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1843_ (.A1(_0558_),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1844_ (.A1(_0697_),
    .A2(_0874_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1845_ (.A1(_0580_),
    .A2(_0814_),
    .B1(_0921_),
    .B2(_0628_),
    .C(_0689_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1846_ (.A1(_0570_),
    .A2(_0761_),
    .B(_0784_),
    .C(_0590_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1847_ (.A1(_0922_),
    .A2(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1848_ (.A1(_0603_),
    .A2(_0606_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1849_ (.I(_0748_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1850_ (.A1(_0925_),
    .A2(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1851_ (.A1(_0866_),
    .A2(_0606_),
    .A3(_0800_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1852_ (.A1(_0815_),
    .A2(_0927_),
    .B(_0928_),
    .C(_0811_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1853_ (.A1(_0772_),
    .A2(_0924_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1854_ (.A1(_0920_),
    .A2(_0930_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1855_ (.A1(_0739_),
    .A2(_0752_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1856_ (.A1(_0881_),
    .A2(_0887_),
    .B(_0806_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1857_ (.I(_0708_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1858_ (.A1(_0932_),
    .A2(_0933_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1859_ (.I(_0885_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1860_ (.A1(_0839_),
    .A2(_0840_),
    .B1(_0926_),
    .B2(_0882_),
    .C(_0849_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1861_ (.A1(_0622_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1862_ (.A1(_0819_),
    .A2(_0824_),
    .B(_0737_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1863_ (.I(_0611_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1864_ (.A1(_0590_),
    .A2(_0685_),
    .A3(_0603_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1865_ (.A1(_0940_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1866_ (.A1(_0759_),
    .A2(_0942_),
    .B(_0716_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1867_ (.A1(_0936_),
    .A2(_0938_),
    .B1(_0939_),
    .B2(_0696_),
    .C(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1868_ (.A1(_0769_),
    .A2(_0818_),
    .A3(_0822_),
    .A4(_0718_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1869_ (.A1(_0849_),
    .A2(_0870_),
    .B(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _1870_ (.A1(_0885_),
    .A2(_0946_),
    .B1(_0802_),
    .B2(_0789_),
    .C1(_0801_),
    .C2(_0591_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1871_ (.A1(_0906_),
    .A2(_0818_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1872_ (.A1(_0882_),
    .A2(_0804_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1873_ (.A1(_0844_),
    .A2(_0741_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _1874_ (.I0(_0908_),
    .I1(_0948_),
    .I2(_0949_),
    .I3(_0950_),
    .S0(_0765_),
    .S1(_0912_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1875_ (.I(_0903_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1876_ (.A1(_0623_),
    .A2(_0673_),
    .A3(_0879_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1877_ (.A1(_0805_),
    .A2(_0947_),
    .B1(_0951_),
    .B2(_0952_),
    .C(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1878_ (.A1(_0556_),
    .A2(_0954_),
    .B(_0944_),
    .C(_0807_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1879_ (.A1(_0542_),
    .A2(_0796_),
    .B1(_0935_),
    .B2(_0944_),
    .C(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1880_ (.A1(_0890_),
    .A2(_0931_),
    .A3(_0956_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1881_ (.A1(_0897_),
    .A2(_0956_),
    .B(_0931_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1882_ (.A1(_0918_),
    .A2(_0957_),
    .A3(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1883_ (.I(_0957_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1884_ (.A1(_0960_),
    .A2(_0958_),
    .B(_0918_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1885_ (.A1(_0877_),
    .A2(_0897_),
    .A3(_0895_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1886_ (.A1(_0863_),
    .A2(_0898_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1887_ (.A1(_0959_),
    .A2(_0961_),
    .A3(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1888_ (.A1(_0959_),
    .A2(_0961_),
    .B(_0963_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1889_ (.A1(_0964_),
    .A2(_0965_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1890_ (.A1(_0863_),
    .A2(_0896_),
    .A3(_0898_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1891_ (.A1(_0896_),
    .A2(_0898_),
    .B(_0863_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1892_ (.A1(_0838_),
    .A2(_0967_),
    .A3(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1893_ (.A1(_0835_),
    .A2(_0900_),
    .B(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1894_ (.A1(_0966_),
    .A2(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1895_ (.I(_0971_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1896_ (.A1(_0918_),
    .A2(_0957_),
    .A3(_0958_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1897_ (.A1(_0960_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1898_ (.A1(_0866_),
    .A2(_0578_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1899_ (.A1(_0570_),
    .A2(_0814_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1900_ (.A1(_0974_),
    .A2(_0867_),
    .A3(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1901_ (.A1(_0734_),
    .A2(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1902_ (.A1(_0588_),
    .A2(_0743_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1903_ (.A1(_0815_),
    .A2(_0907_),
    .B(_0767_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1904_ (.A1(_0842_),
    .A2(_0824_),
    .B1(_0978_),
    .B2(_0979_),
    .C(_0772_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1905_ (.A1(_0977_),
    .A2(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1906_ (.A1(_0919_),
    .A2(_0930_),
    .B(_0558_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1907_ (.A1(_0981_),
    .A2(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1908_ (.A1(_0557_),
    .A2(_0954_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(_0668_),
    .A2(_0742_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1910_ (.A1(_0577_),
    .A2(_0700_),
    .B(_0697_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1911_ (.A1(_0941_),
    .A2(_0986_),
    .B(_0587_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1912_ (.A1(_0720_),
    .A2(_0735_),
    .A3(_0781_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1913_ (.A1(_0596_),
    .A2(_0631_),
    .A3(_0907_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1914_ (.A1(_0988_),
    .A2(_0989_),
    .B(_0593_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1915_ (.A1(_0613_),
    .A2(_0988_),
    .A3(_0989_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1916_ (.A1(_0987_),
    .A2(_0990_),
    .B(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1917_ (.A1(_0811_),
    .A2(_0985_),
    .B1(_0992_),
    .B2(_0885_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1918_ (.A1(_0934_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1919_ (.A1(_0984_),
    .A2(_0993_),
    .B(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1920_ (.A1(_0891_),
    .A2(_0894_),
    .B(_0655_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1921_ (.A1(_0892_),
    .A2(_0995_),
    .B(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1922_ (.I(_0757_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1923_ (.A1(_0852_),
    .A2(_0857_),
    .A3(_0860_),
    .A4(_0916_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1924_ (.A1(_0998_),
    .A2(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1925_ (.I(_0866_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1926_ (.A1(_1001_),
    .A2(_0692_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1927_ (.A1(_0940_),
    .A2(_0925_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1928_ (.A1(_1002_),
    .A2(_1003_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1929_ (.I(_0614_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1930_ (.A1(_0729_),
    .A2(_0743_),
    .B(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1931_ (.I(_0725_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1932_ (.A1(_0571_),
    .A2(_0907_),
    .A3(_0718_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1933_ (.A1(_1007_),
    .A2(_0728_),
    .B1(_1008_),
    .B2(_0882_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1934_ (.A1(_0712_),
    .A2(_1006_),
    .B1(_1009_),
    .B2(_1005_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1935_ (.A1(_0812_),
    .A2(_1004_),
    .B1(_1010_),
    .B2(_0936_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1936_ (.A1(_0998_),
    .A2(_0999_),
    .A3(_1011_),
    .B(\p_shaping_Q.p_shaping_I.counter[1] ),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1937_ (.A1(_1000_),
    .A2(_1011_),
    .B(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1938_ (.A1(_0983_),
    .A2(_0997_),
    .A3(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1939_ (.A1(_0973_),
    .A2(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1940_ (.A1(_0959_),
    .A2(_0961_),
    .A3(_0963_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1941_ (.A1(_0966_),
    .A2(_0970_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1942_ (.A1(_1016_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1943_ (.A1(_1015_),
    .A2(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1944_ (.I(_1019_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1945_ (.A1(_0933_),
    .A2(_0993_),
    .B(_0708_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1946_ (.A1(_0839_),
    .A2(_0671_),
    .B(_0908_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1947_ (.A1(_0600_),
    .A2(_0840_),
    .B(_0812_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1948_ (.A1(_0765_),
    .A2(_0614_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1949_ (.A1(_0906_),
    .A2(_0659_),
    .A3(_0825_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1950_ (.A1(_0825_),
    .A2(_0759_),
    .B(_0748_),
    .C(_0613_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1951_ (.A1(_1024_),
    .A2(_1025_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1952_ (.A1(_0661_),
    .A2(_1023_),
    .B(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1953_ (.A1(_1021_),
    .A2(_1022_),
    .B1(_1027_),
    .B2(_0851_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1954_ (.A1(_1020_),
    .A2(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1955_ (.A1(_0892_),
    .A2(_1029_),
    .B(_0996_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1956_ (.A1(_0919_),
    .A2(_0930_),
    .A3(_0977_),
    .A4(_0980_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1957_ (.A1(_0704_),
    .A2(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1958_ (.A1(_0853_),
    .A2(_1007_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1959_ (.I(_0537_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1960_ (.A1(_1001_),
    .A2(_0599_),
    .B1(_1033_),
    .B2(_1034_),
    .C(_0912_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1961_ (.A1(_0849_),
    .A2(_0515_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1962_ (.A1(_0912_),
    .A2(_0903_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1963_ (.A1(_0851_),
    .A2(_1035_),
    .A3(_1036_),
    .B1(_1037_),
    .B2(_0987_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1964_ (.I0(_1032_),
    .I1(_0559_),
    .S(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1965_ (.A1(_1030_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1966_ (.A1(_0999_),
    .A2(_1011_),
    .B(_0757_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1967_ (.I(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1968_ (.I(_1002_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1969_ (.I(_0940_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1970_ (.I(_0853_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1971_ (.A1(_1045_),
    .A2(_0913_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1972_ (.A1(_1044_),
    .A2(_0948_),
    .A3(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1973_ (.I(_1005_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1974_ (.A1(_1048_),
    .A2(_0874_),
    .A3(_0926_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1975_ (.A1(_1047_),
    .A2(_1049_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1976_ (.I(_1048_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1977_ (.A1(_1051_),
    .A2(_0762_),
    .B1(_1047_),
    .B2(_1049_),
    .C(_0936_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1978_ (.A1(_1043_),
    .A2(_1037_),
    .B1(_1050_),
    .B2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1979_ (.A1(_1041_),
    .A2(_1053_),
    .B(_0566_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1980_ (.A1(_1042_),
    .A2(_1053_),
    .B(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1981_ (.A1(_1040_),
    .A2(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1982_ (.A1(_0983_),
    .A2(_0997_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1983_ (.I(_1013_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1984_ (.A1(_0983_),
    .A2(_0997_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1985_ (.A1(_1057_),
    .A2(_1058_),
    .B(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1986_ (.A1(_1056_),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1987_ (.A1(_0960_),
    .A2(_0972_),
    .B(_1014_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1988_ (.A1(_0960_),
    .A2(_0972_),
    .A3(_1014_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1989_ (.A1(_1016_),
    .A2(_1017_),
    .A3(_1062_),
    .B(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1990_ (.A1(_1061_),
    .A2(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1991_ (.I(_1065_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1992_ (.A1(_0864_),
    .A2(_1031_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1993_ (.I(_0851_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1994_ (.A1(_1005_),
    .A2(_0870_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1995_ (.A1(_1043_),
    .A2(_0826_),
    .B(_0762_),
    .C(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1996_ (.A1(_0952_),
    .A2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1997_ (.I(_0539_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1998_ (.A1(_1067_),
    .A2(_0926_),
    .B(_1070_),
    .C(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1999_ (.A1(_1066_),
    .A2(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2000_ (.I(_1020_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2001_ (.I(_0842_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2002_ (.A1(_0769_),
    .A2(_0867_),
    .A3(_0904_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2003_ (.A1(_0940_),
    .A2(_0847_),
    .B(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2004_ (.I(_0921_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2005_ (.A1(_0571_),
    .A2(_0665_),
    .B1(_0904_),
    .B2(_1078_),
    .C(_0842_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2006_ (.A1(_1075_),
    .A2(_1077_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2007_ (.A1(_0936_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2008_ (.A1(_0819_),
    .A2(_0588_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2009_ (.A1(_0952_),
    .A2(_1068_),
    .A3(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2010_ (.A1(_1081_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2011_ (.I0(_1074_),
    .I1(_0934_),
    .S(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2012_ (.A1(_0806_),
    .A2(_0807_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2013_ (.A1(_0797_),
    .A2(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2014_ (.A1(_0655_),
    .A2(_1087_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2015_ (.A1(_0892_),
    .A2(_1085_),
    .B(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2016_ (.I(_1067_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2017_ (.A1(_1075_),
    .A2(_0628_),
    .A3(_1046_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2018_ (.I(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2019_ (.A1(_0905_),
    .A2(_1036_),
    .B1(_1092_),
    .B2(_1078_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2020_ (.A1(_1090_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2021_ (.A1(_1041_),
    .A2(_1094_),
    .B(_0566_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2022_ (.A1(_1042_),
    .A2(_1094_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2023_ (.A1(_1073_),
    .A2(_1089_),
    .A3(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2024_ (.A1(_1030_),
    .A2(_1039_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2025_ (.A1(_1040_),
    .A2(_1055_),
    .B(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2026_ (.A1(_1097_),
    .A2(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2027_ (.A1(_1056_),
    .A2(_1060_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2028_ (.A1(_1061_),
    .A2(_1064_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2029_ (.A1(_1101_),
    .A2(_1102_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2030_ (.A1(_1100_),
    .A2(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2031_ (.I(_1104_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2032_ (.A1(_0819_),
    .A2(_0712_),
    .B1(_0927_),
    .B2(_1044_),
    .C(_1075_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2033_ (.A1(_1031_),
    .A2(_1105_),
    .B(_0864_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2034_ (.I0(_0864_),
    .I1(_1106_),
    .S(_0540_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2035_ (.A1(_0622_),
    .A2(_1076_),
    .B(_0952_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2036_ (.A1(_0668_),
    .A2(_0716_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2037_ (.A1(_0844_),
    .A2(_0696_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2038_ (.A1(_1001_),
    .A2(_0662_),
    .B(_0746_),
    .C(_0728_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2039_ (.A1(_0847_),
    .A2(_1109_),
    .B1(_0986_),
    .B2(_1110_),
    .C(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2040_ (.A1(_1108_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2041_ (.I0(_0934_),
    .I1(_1074_),
    .S(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2042_ (.A1(_0893_),
    .A2(_1114_),
    .B(_0996_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2043_ (.A1(_1107_),
    .A2(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2044_ (.I(_1090_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2045_ (.A1(_1001_),
    .A2(_0840_),
    .B(_0974_),
    .C(_1051_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2046_ (.I(_1075_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2047_ (.A1(_0607_),
    .A2(_1078_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2048_ (.A1(_0999_),
    .A2(_1011_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2049_ (.A1(_0938_),
    .A2(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2050_ (.A1(_1117_),
    .A2(_1118_),
    .A3(_1120_),
    .B1(_1122_),
    .B2(_0998_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2051_ (.A1(_1090_),
    .A2(_0998_),
    .A3(_1118_),
    .A4(_1120_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2052_ (.A1(_0756_),
    .A2(_1123_),
    .A3(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2053_ (.A1(_1116_),
    .A2(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2054_ (.A1(_1073_),
    .A2(_1089_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2055_ (.A1(_1073_),
    .A2(_1089_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2056_ (.A1(_1127_),
    .A2(_1128_),
    .A3(_1096_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2057_ (.A1(_1127_),
    .A2(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2058_ (.A1(_1126_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2059_ (.A1(_1040_),
    .A2(_1055_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2060_ (.A1(_1098_),
    .A2(_1132_),
    .A3(_1097_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2061_ (.A1(_1061_),
    .A2(_1100_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2062_ (.A1(_1016_),
    .A2(_1062_),
    .B(_1063_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2063_ (.A1(_0966_),
    .A2(_0970_),
    .A3(_1015_),
    .B(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2064_ (.A1(_1098_),
    .A2(_1132_),
    .B(_1097_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2065_ (.A1(_1101_),
    .A2(_1133_),
    .B1(_1134_),
    .B2(_1136_),
    .C(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2066_ (.A1(_1131_),
    .A2(_1138_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2067_ (.I(_1139_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2068_ (.I(_1115_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2069_ (.A1(_1107_),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2070_ (.A1(_1116_),
    .A2(_1125_),
    .B(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2071_ (.I(_1067_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2072_ (.A1(_1143_),
    .A2(_0677_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2073_ (.I(_1044_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2074_ (.A1(_1145_),
    .A2(_1045_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2075_ (.A1(_1143_),
    .A2(_1146_),
    .A3(_1043_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2076_ (.A1(_1071_),
    .A2(_1144_),
    .A3(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2077_ (.I0(_0559_),
    .I1(_1032_),
    .S(_1148_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2078_ (.A1(_1045_),
    .A2(_1007_),
    .B(_0728_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2079_ (.A1(_1048_),
    .A2(_0729_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2080_ (.A1(_1048_),
    .A2(_0607_),
    .B1(_1150_),
    .B2(_1151_),
    .C(_1067_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2081_ (.A1(_1143_),
    .A2(_1105_),
    .B(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2082_ (.A1(_1074_),
    .A2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2083_ (.A1(_0557_),
    .A2(_1153_),
    .B(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2084_ (.A1(_0893_),
    .A2(_1155_),
    .B(_0996_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2085_ (.A1(_1149_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2086_ (.I(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2087_ (.A1(_0638_),
    .A2(_0740_),
    .B(_0824_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2088_ (.A1(_1119_),
    .A2(_1078_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2089_ (.A1(_1119_),
    .A2(_1159_),
    .B(_1160_),
    .C(_1117_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2090_ (.A1(_1042_),
    .A2(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2091_ (.A1(_0859_),
    .A2(_1161_),
    .B(_1162_),
    .C(_0567_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2092_ (.A1(_1158_),
    .A2(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2093_ (.A1(_1142_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2094_ (.A1(_1142_),
    .A2(_1164_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2095_ (.A1(_1165_),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2096_ (.A1(_1126_),
    .A2(_1130_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2097_ (.A1(_1131_),
    .A2(_1138_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2098_ (.A1(_1168_),
    .A2(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2099_ (.A1(_1167_),
    .A2(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2100_ (.I(_1171_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2101_ (.A1(_1071_),
    .A2(_1066_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2102_ (.A1(_0559_),
    .A2(_1071_),
    .B1(_0677_),
    .B2(_1117_),
    .C(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2103_ (.A1(_1043_),
    .A2(_1003_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2104_ (.A1(_1044_),
    .A2(_0826_),
    .B(_1036_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2105_ (.A1(_0713_),
    .A2(_1174_),
    .B1(_1175_),
    .B2(_1143_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2106_ (.A1(_0797_),
    .A2(_1020_),
    .B(_1087_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2107_ (.A1(_1176_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2108_ (.A1(_0007_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2109_ (.A1(_1173_),
    .A2(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2110_ (.A1(_1051_),
    .A2(_0621_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2111_ (.A1(_1090_),
    .A2(_1160_),
    .A3(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2112_ (.A1(_1042_),
    .A2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2113_ (.A1(_0859_),
    .A2(_1182_),
    .B(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2114_ (.A1(_0756_),
    .A2(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2115_ (.I(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2116_ (.A1(_1180_),
    .A2(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2117_ (.A1(_1158_),
    .A2(_1163_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2118_ (.A1(_1149_),
    .A2(_1156_),
    .B(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2119_ (.A1(_1187_),
    .A2(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2120_ (.I(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2121_ (.A1(_1126_),
    .A2(_1130_),
    .B(_1165_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2122_ (.A1(_1169_),
    .A2(_1192_),
    .B(_1166_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2123_ (.A1(_1191_),
    .A2(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2124_ (.I(_1194_),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2125_ (.I(_1173_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2126_ (.A1(_1195_),
    .A2(_1179_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2127_ (.A1(_1180_),
    .A2(_1186_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2128_ (.A1(_0713_),
    .A2(_1003_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2129_ (.A1(_0617_),
    .A2(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2130_ (.A1(_1074_),
    .A2(_1199_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2131_ (.A1(_0557_),
    .A2(_1199_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2132_ (.A1(_0893_),
    .A2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2133_ (.A1(_1201_),
    .A2(_1203_),
    .B(_0897_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2134_ (.A1(_1195_),
    .A2(_1185_),
    .A3(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2135_ (.A1(_1196_),
    .A2(_1197_),
    .B(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2136_ (.A1(_1196_),
    .A2(_1197_),
    .A3(_1205_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2137_ (.A1(_1206_),
    .A2(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2138_ (.A1(_1187_),
    .A2(_1189_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2139_ (.A1(_1191_),
    .A2(_1193_),
    .B(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2140_ (.A1(_1208_),
    .A2(_1210_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2141_ (.I(_1212_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2142_ (.A1(_1186_),
    .A2(_1204_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2143_ (.A1(_1186_),
    .A2(_1204_),
    .B(_1195_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2144_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2145_ (.A1(_1196_),
    .A2(_1197_),
    .A3(_1205_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2146_ (.A1(_1190_),
    .A2(_1208_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2147_ (.A1(_1209_),
    .A2(_1216_),
    .B1(_1217_),
    .B2(_1193_),
    .C(_1206_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2148_ (.A1(_0656_),
    .A2(_1177_),
    .B1(_1215_),
    .B2(_1218_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2149_ (.A1(_0684_),
    .A2(_0777_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2150_ (.I(_1219_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2151_ (.I(net32),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2152_ (.A1(_1221_),
    .A2(_0140_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2153_ (.I(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2154_ (.A1(_1296_),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2155_ (.A1(_1350_),
    .A2(_1372_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2156_ (.I(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2157_ (.A1(_1224_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2158_ (.I(net35),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2159_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2160_ (.I(_1229_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2161_ (.I(_0140_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2162_ (.I(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2163_ (.A1(_0129_),
    .A2(_1372_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2164_ (.I(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2165_ (.A1(_1233_),
    .A2(_1235_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2166_ (.I(_1361_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2167_ (.I(_0270_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2168_ (.I(_1307_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2169_ (.A1(_1237_),
    .A2(_1238_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2170_ (.I(_0205_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2171_ (.A1(_1231_),
    .A2(_1236_),
    .A3(_1240_),
    .B(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2172_ (.I(_1339_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2173_ (.I(_1350_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2174_ (.I(net34),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2175_ (.A1(_1245_),
    .A2(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2176_ (.I(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2177_ (.I(_1285_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2178_ (.A1(_1249_),
    .A2(_1222_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2179_ (.I(_1245_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2180_ (.I(_1221_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2181_ (.A1(_1251_),
    .A2(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2182_ (.A1(_1244_),
    .A2(_1248_),
    .B(_1250_),
    .C(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2183_ (.I(_1242_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2184_ (.I(net53),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2185_ (.I(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2186_ (.I(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2187_ (.A1(_1227_),
    .A2(_1243_),
    .B1(_1255_),
    .B2(_1256_),
    .C(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2188_ (.I(_0129_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2189_ (.A1(_1261_),
    .A2(_1211_),
    .A3(_1232_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2190_ (.I(_0259_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2191_ (.I(_1232_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2192_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2193_ (.A1(_1264_),
    .A2(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2194_ (.I(_1285_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2195_ (.I(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2196_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2197_ (.A1(_1267_),
    .A2(_0162_),
    .B(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2198_ (.A1(_1245_),
    .A2(_1221_),
    .A3(_1246_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2199_ (.I(net36),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2200_ (.A1(_1228_),
    .A2(_1272_),
    .B(_1273_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2201_ (.A1(_0216_),
    .A2(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2202_ (.A1(_1262_),
    .A2(_1271_),
    .B(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2203_ (.A1(_1260_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2204_ (.A1(\p_shaping_I.p_shaping_I.counter[1] ),
    .A2(\p_shaping_I.p_shaping_I.counter[0] ),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2205_ (.I(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2206_ (.I(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2207_ (.A1(_1278_),
    .A2(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2208_ (.A1(_0118_),
    .A2(_0183_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2209_ (.I(_1234_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2210_ (.A1(_1318_),
    .A2(_1284_),
    .B(_1339_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2211_ (.I(_1252_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2212_ (.A1(_1350_),
    .A2(net32),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2213_ (.I(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2214_ (.A1(_1287_),
    .A2(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2215_ (.I(_1273_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2216_ (.I(_1241_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2217_ (.A1(_1237_),
    .A2(_1268_),
    .A3(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2218_ (.A1(_1286_),
    .A2(_1290_),
    .B(_1291_),
    .C(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2219_ (.I(_1211_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2220_ (.A1(_1361_),
    .A2(_1253_),
    .B(_1232_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2221_ (.A1(_1295_),
    .A2(_1297_),
    .B(_0205_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2222_ (.A1(_1258_),
    .A2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2223_ (.I(_0032_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2224_ (.A1(_1300_),
    .A2(_1287_),
    .B(_1295_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2225_ (.I0(_1221_),
    .I1(_0129_),
    .S(_0140_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2226_ (.I(_1302_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2227_ (.A1(_1229_),
    .A2(_1284_),
    .A3(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2228_ (.A1(_1240_),
    .A2(_1301_),
    .B(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2229_ (.A1(_1283_),
    .A2(_1294_),
    .B1(_1299_),
    .B2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2230_ (.I(\p_shaping_I.p_shaping_I.counter[1] ),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2231_ (.A1(_1249_),
    .A2(_1225_),
    .B(_0087_),
    .C(_1252_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2232_ (.A1(_1245_),
    .A2(_0032_),
    .B(_1285_),
    .C(_1246_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2233_ (.A1(_0076_),
    .A2(_1310_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2234_ (.I(_1200_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2235_ (.A1(_0281_),
    .A2(_1312_),
    .A3(_1247_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2236_ (.A1(_0173_),
    .A2(_1262_),
    .A3(_1309_),
    .B1(_1311_),
    .B2(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2237_ (.I(_1211_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2238_ (.A1(_1312_),
    .A2(_0076_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2239_ (.A1(_1315_),
    .A2(_1254_),
    .B1(_1316_),
    .B2(_0216_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2240_ (.A1(_1314_),
    .A2(_1317_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2241_ (.A1(_1308_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2242_ (.A1(_1306_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2243_ (.A1(_1282_),
    .A2(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2244_ (.I(_1322_),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2245_ (.I(_0087_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2246_ (.I(_1323_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2247_ (.I(_1291_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2248_ (.A1(_1266_),
    .A2(_1226_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2249_ (.A1(_0259_),
    .A2(_0291_),
    .A3(_1263_),
    .B(_1315_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2250_ (.I(_0032_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2251_ (.A1(_1237_),
    .A2(_1329_),
    .B(_1318_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2252_ (.A1(_1269_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2253_ (.A1(_1327_),
    .A2(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2254_ (.A1(_1325_),
    .A2(_1326_),
    .A3(_1332_),
    .B(_0183_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2255_ (.I(_1261_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2256_ (.I(_1329_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2257_ (.A1(_1334_),
    .A2(_1335_),
    .A3(_1266_),
    .B(_1250_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2258_ (.I(_1268_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2259_ (.I(_1246_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2260_ (.A1(_1251_),
    .A2(_1338_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2261_ (.A1(_1335_),
    .A2(_1337_),
    .A3(_1340_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2262_ (.A1(_1336_),
    .A2(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2263_ (.A1(_1273_),
    .A2(_0087_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2264_ (.I(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2265_ (.I(_1239_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2266_ (.A1(_1334_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2267_ (.I(_0043_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2268_ (.A1(_1231_),
    .A2(_1347_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2269_ (.A1(_1270_),
    .A2(_1346_),
    .B(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2270_ (.I(_0227_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2271_ (.A1(_1324_),
    .A2(_1333_),
    .B1(_1342_),
    .B2(_1344_),
    .C1(_1349_),
    .C2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2272_ (.A1(_1260_),
    .A2(_1277_),
    .B(net44),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2273_ (.A1(_1352_),
    .A2(_1353_),
    .B(_1280_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2274_ (.A1(_1352_),
    .A2(_1353_),
    .B(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2275_ (.A1(_1228_),
    .A2(_1252_),
    .A3(_1288_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2276_ (.A1(_1312_),
    .A2(_1302_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2277_ (.A1(_1310_),
    .A2(_1356_),
    .A3(_1357_),
    .B(_1323_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2278_ (.I(_1261_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2279_ (.I(_1253_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2280_ (.A1(_1359_),
    .A2(_1360_),
    .B(_1315_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2281_ (.I(_1228_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2282_ (.A1(_1363_),
    .A2(_1347_),
    .B(_0216_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2283_ (.A1(_1362_),
    .A2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2284_ (.A1(_1358_),
    .A2(_1365_),
    .B(_1325_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2285_ (.A1(_1269_),
    .A2(_0162_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2286_ (.A1(_1300_),
    .A2(_1265_),
    .B(_1359_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2287_ (.A1(_1244_),
    .A2(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2288_ (.A1(_0173_),
    .A2(_1257_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2289_ (.I(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2290_ (.A1(_1367_),
    .A2(_1369_),
    .B(_1371_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2291_ (.A1(_1366_),
    .A2(_0022_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2292_ (.A1(_0552_),
    .A2(_1306_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2293_ (.A1(_0023_),
    .A2(_0024_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2294_ (.I(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2295_ (.A1(_1314_),
    .A2(_1317_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2296_ (.I(_1261_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2297_ (.A1(_0028_),
    .A2(_1249_),
    .A3(_1338_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2298_ (.A1(_1251_),
    .A2(_0281_),
    .B(_1312_),
    .C(_1292_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2299_ (.A1(_1360_),
    .A2(_0029_),
    .B(_0030_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2300_ (.A1(_0173_),
    .A2(_1356_),
    .A3(_1357_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2301_ (.A1(_1339_),
    .A2(_0076_),
    .A3(_1289_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2302_ (.A1(_0118_),
    .A2(_0034_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2303_ (.A1(_1276_),
    .A2(_0031_),
    .B1(_0033_),
    .B2(_0035_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2304_ (.A1(_0026_),
    .A2(_0027_),
    .B(_0036_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2305_ (.A1(_0026_),
    .A2(_0027_),
    .A3(_0036_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2306_ (.A1(_1308_),
    .A2(_0037_),
    .A3(_0038_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2307_ (.A1(_1355_),
    .A2(_0025_),
    .A3(_0039_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2308_ (.I(_1308_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2309_ (.A1(_0041_),
    .A2(_1306_),
    .A3(_1319_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2310_ (.A1(_1282_),
    .A2(_1321_),
    .B(_0042_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2311_ (.A1(_0040_),
    .A2(_0044_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2312_ (.A1(_0025_),
    .A2(_0039_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2313_ (.A1(_0025_),
    .A2(_0039_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2314_ (.A1(_1355_),
    .A2(_0046_),
    .B(_0047_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2315_ (.A1(_0544_),
    .A2(_0553_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2316_ (.A1(_0324_),
    .A2(_0049_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2317_ (.I(_1273_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2318_ (.A1(_1292_),
    .A2(_1225_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2319_ (.A1(_1238_),
    .A2(_1239_),
    .B(_1295_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2320_ (.A1(_0052_),
    .A2(_0053_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2321_ (.I(_0281_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2322_ (.A1(_1251_),
    .A2(_1338_),
    .B(_1249_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2323_ (.A1(_0205_),
    .A2(_0057_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2324_ (.A1(_1363_),
    .A2(_1248_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2325_ (.A1(_0056_),
    .A2(_0058_),
    .A3(_0059_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2326_ (.A1(_0051_),
    .A2(_0055_),
    .B(_0060_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2327_ (.A1(_1244_),
    .A2(_0227_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2328_ (.A1(_1238_),
    .A2(_1263_),
    .B(_1237_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2329_ (.A1(_1292_),
    .A2(_1288_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2330_ (.A1(_1220_),
    .A2(_0064_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2331_ (.A1(_0028_),
    .A2(_1329_),
    .A3(_1295_),
    .A4(_1287_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2332_ (.A1(_1291_),
    .A2(_0067_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2333_ (.A1(_0066_),
    .A2(_0068_),
    .B(_1259_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2334_ (.A1(_1259_),
    .A2(_0061_),
    .B1(_0062_),
    .B2(_0063_),
    .C(_0069_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2335_ (.A1(_1278_),
    .A2(_1352_),
    .B(_0548_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2336_ (.A1(_0050_),
    .A2(_0070_),
    .A3(_0071_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2337_ (.A1(_1306_),
    .A2(_1366_),
    .A3(_0022_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2338_ (.A1(_0545_),
    .A2(_0073_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2339_ (.I(_1290_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2340_ (.A1(_1370_),
    .A2(_1286_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2341_ (.A1(_1318_),
    .A2(_1284_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2342_ (.A1(_1327_),
    .A2(_0078_),
    .B(_1364_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2343_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2344_ (.A1(_1238_),
    .A2(_1247_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2345_ (.A1(_1300_),
    .A2(_1229_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2346_ (.A1(_1337_),
    .A2(_0080_),
    .B1(_0081_),
    .B2(_0082_),
    .C(_0118_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2347_ (.A1(_0079_),
    .A2(_0083_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2348_ (.A1(_0075_),
    .A2(_0077_),
    .B1(_0084_),
    .B2(_1242_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2349_ (.I(_0085_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2350_ (.I(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2351_ (.A1(_1307_),
    .A2(_1234_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2352_ (.A1(_1220_),
    .A2(_0078_),
    .B1(_0089_),
    .B2(_0030_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2353_ (.A1(_0028_),
    .A2(_1329_),
    .B(_1287_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2354_ (.A1(_1220_),
    .A2(_0091_),
    .B(_1250_),
    .C(_1291_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2355_ (.A1(_1268_),
    .A2(_1284_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2356_ (.A1(_0028_),
    .A2(_1253_),
    .B(_1338_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2357_ (.A1(_1223_),
    .A2(_0093_),
    .B1(_0094_),
    .B2(_1224_),
    .C(_1343_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2358_ (.A1(_1370_),
    .A2(_0090_),
    .B1(_0092_),
    .B2(_1258_),
    .C(_0095_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2359_ (.A1(_1314_),
    .A2(_1317_),
    .B1(_0033_),
    .B2(_0035_),
    .C1(_0031_),
    .C2(_1276_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2360_ (.A1(_0088_),
    .A2(_0096_),
    .A3(_0097_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2361_ (.A1(_0088_),
    .A2(_0097_),
    .B(_0096_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2362_ (.A1(\p_shaping_I.p_shaping_I.counter[1] ),
    .A2(_0099_),
    .A3(_0100_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2363_ (.A1(_0074_),
    .A2(_0086_),
    .A3(_0101_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2364_ (.A1(_1281_),
    .A2(_0072_),
    .A3(_0102_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2365_ (.I(_1281_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2366_ (.A1(_0021_),
    .A2(_0072_),
    .B(_0102_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2367_ (.A1(_0103_),
    .A2(_0104_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2368_ (.A1(_0045_),
    .A2(_0048_),
    .A3(_0105_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2369_ (.I(_0106_),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2370_ (.A1(_0103_),
    .A2(_0104_),
    .B(_0048_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2371_ (.A1(_0048_),
    .A2(_0103_),
    .A3(_0104_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2372_ (.A1(_0045_),
    .A2(_0108_),
    .B(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2373_ (.A1(_0074_),
    .A2(_0086_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2374_ (.A1(_0111_),
    .A2(_0101_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2375_ (.A1(_0112_),
    .A2(_0103_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2376_ (.I(_0070_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2377_ (.A1(_1278_),
    .A2(_1352_),
    .A3(_0114_),
    .B(_0548_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2378_ (.A1(_1324_),
    .A2(_1275_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2379_ (.I(_1326_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2380_ (.A1(_0117_),
    .A2(_1331_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2381_ (.I(_1325_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2382_ (.A1(_0120_),
    .A2(_1346_),
    .A3(_1293_),
    .A4(_0052_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2383_ (.I(_1259_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2384_ (.A1(_1270_),
    .A2(_1223_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2385_ (.A1(_1313_),
    .A2(_0123_),
    .B(_0120_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2386_ (.A1(_0122_),
    .A2(_0124_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2387_ (.A1(_0116_),
    .A2(_1293_),
    .A3(_0119_),
    .B1(_0121_),
    .B2(_0125_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2388_ (.A1(_0115_),
    .A2(_0126_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2389_ (.A1(_0050_),
    .A2(_0127_),
    .B(_1281_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2390_ (.A1(net46),
    .A2(_0049_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2391_ (.A1(_0115_),
    .A2(_0126_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2392_ (.A1(_0130_),
    .A2(_0131_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2393_ (.A1(_0128_),
    .A2(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2394_ (.A1(_1360_),
    .A2(_1248_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2395_ (.A1(_1269_),
    .A2(_1235_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2396_ (.A1(_1345_),
    .A2(_0302_),
    .A3(_1362_),
    .B1(_0134_),
    .B2(_0135_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2397_ (.A1(_1325_),
    .A2(_0136_),
    .B(_0067_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2398_ (.I(_1363_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2399_ (.A1(_1359_),
    .A2(_1300_),
    .B(_1239_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2400_ (.I(_0081_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2401_ (.A1(_1231_),
    .A2(_0141_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2402_ (.A1(_0138_),
    .A2(_0139_),
    .B(_0142_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2403_ (.A1(_0291_),
    .A2(_1233_),
    .B(_1315_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2404_ (.A1(_1335_),
    .A2(_0029_),
    .B1(_0144_),
    .B2(_1254_),
    .C(_1272_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2405_ (.A1(_1323_),
    .A2(_0137_),
    .B1(_0143_),
    .B2(_1343_),
    .C1(_0145_),
    .C2(_1351_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2406_ (.A1(_0073_),
    .A2(_0086_),
    .B(_0546_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2407_ (.A1(_0146_),
    .A2(_0147_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2408_ (.A1(_0051_),
    .A2(_1258_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2409_ (.A1(_1265_),
    .A2(_1226_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2410_ (.A1(_0056_),
    .A2(_1233_),
    .B1(_0063_),
    .B2(_1337_),
    .C(_0150_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2411_ (.A1(_0056_),
    .A2(_1233_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2412_ (.I(_0064_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2413_ (.A1(_0153_),
    .A2(_0154_),
    .B(_1368_),
    .C(_1244_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2414_ (.A1(_0149_),
    .A2(_0152_),
    .A3(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2415_ (.A1(_0259_),
    .A2(_1263_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2416_ (.A1(_1337_),
    .A2(_0157_),
    .A3(_0139_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2417_ (.A1(_0291_),
    .A2(_1265_),
    .B(_1229_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2418_ (.A1(_0162_),
    .A2(_0159_),
    .B(_1370_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2419_ (.A1(_1286_),
    .A2(_1290_),
    .A3(_1303_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2420_ (.A1(_1363_),
    .A2(_1303_),
    .B(_1343_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2421_ (.I(_0163_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2422_ (.A1(_0158_),
    .A2(_0160_),
    .B1(_0161_),
    .B2(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2423_ (.A1(_0156_),
    .A2(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2424_ (.A1(_0096_),
    .A2(_0097_),
    .B(_0088_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2425_ (.A1(_0166_),
    .A2(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2426_ (.A1(_1308_),
    .A2(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2427_ (.A1(_0148_),
    .A2(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2428_ (.A1(_0113_),
    .A2(_0133_),
    .A3(_0170_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2429_ (.A1(_0110_),
    .A2(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2430_ (.I(_0172_),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2431_ (.I(_1256_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2432_ (.A1(_1286_),
    .A2(_0075_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2433_ (.A1(_1345_),
    .A2(_1254_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2434_ (.A1(_0174_),
    .A2(_0157_),
    .A3(_0175_),
    .A4(_0176_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(_1275_),
    .A2(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2436_ (.I(_1230_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2437_ (.I(_1345_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2438_ (.A1(_1230_),
    .A2(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2439_ (.I(_0181_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2440_ (.I(_1264_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2441_ (.A1(_0179_),
    .A2(_0157_),
    .B1(_0182_),
    .B2(_0184_),
    .C(_1344_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2442_ (.A1(_0082_),
    .A2(_1346_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2443_ (.A1(_1351_),
    .A2(_0080_),
    .A3(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2444_ (.A1(_0122_),
    .A2(_0178_),
    .B(_0185_),
    .C(_0187_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2445_ (.A1(_0114_),
    .A2(_0126_),
    .B(_0549_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2446_ (.A1(_0071_),
    .A2(_0189_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2447_ (.A1(_0188_),
    .A2(_0190_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2448_ (.A1(_0130_),
    .A2(_0131_),
    .B(_1279_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2449_ (.A1(_0130_),
    .A2(_0191_),
    .B(_0192_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2450_ (.A1(_0073_),
    .A2(_0085_),
    .A3(_0146_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2451_ (.A1(_0544_),
    .A2(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2452_ (.I(_0029_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2453_ (.I(_1335_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2454_ (.A1(_0180_),
    .A2(_1235_),
    .B1(_0302_),
    .B2(_1301_),
    .C1(_0197_),
    .C2(_0198_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2455_ (.A1(_0051_),
    .A2(_0057_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2456_ (.A1(_0184_),
    .A2(_0200_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2457_ (.I(_1231_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2458_ (.I(_1223_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2459_ (.A1(_1264_),
    .A2(_1274_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2460_ (.A1(_0138_),
    .A2(_1272_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2461_ (.I(_0051_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2462_ (.A1(_0202_),
    .A2(_0203_),
    .B1(_0204_),
    .B2(_0206_),
    .C(_0207_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2463_ (.A1(_0201_),
    .A2(_0208_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2464_ (.A1(_0149_),
    .A2(_0199_),
    .B1(_0209_),
    .B2(_0122_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2465_ (.A1(_0196_),
    .A2(_0210_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2466_ (.I(\p_shaping_I.p_shaping_I.counter[1] ),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2467_ (.A1(_0096_),
    .A2(_0097_),
    .A3(_0156_),
    .A4(_0165_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2468_ (.A1(_0088_),
    .A2(_0213_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2469_ (.A1(_1367_),
    .A2(_0141_),
    .B1(_0052_),
    .B2(_0053_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2470_ (.A1(_0135_),
    .A2(_0200_),
    .B1(_0215_),
    .B2(_0207_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2471_ (.A1(_0138_),
    .A2(_0075_),
    .A3(_0176_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2472_ (.A1(_1256_),
    .A2(_0066_),
    .A3(_0218_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2473_ (.I0(_0217_),
    .I1(_0219_),
    .S(_1323_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2474_ (.A1(_0214_),
    .A2(_0220_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2475_ (.A1(_0212_),
    .A2(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2476_ (.A1(_0211_),
    .A2(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2477_ (.A1(_0193_),
    .A2(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2478_ (.A1(_0148_),
    .A2(_0169_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2479_ (.I(_0128_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2480_ (.A1(_0226_),
    .A2(_0132_),
    .A3(_0170_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2481_ (.A1(_0225_),
    .A2(_0228_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2482_ (.A1(_0224_),
    .A2(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2483_ (.A1(_0226_),
    .A2(_0132_),
    .B(_0170_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2484_ (.A1(_0113_),
    .A2(_0228_),
    .A3(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2485_ (.A1(_0110_),
    .A2(_0171_),
    .B(_0232_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2486_ (.A1(_0230_),
    .A2(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2487_ (.I(_0234_),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2488_ (.A1(_0211_),
    .A2(_0222_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2489_ (.A1(_0193_),
    .A2(_0223_),
    .B(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2490_ (.I(_0050_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2491_ (.I(_0056_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2492_ (.I(_0098_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2493_ (.A1(_0239_),
    .A2(_0181_),
    .B(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2494_ (.A1(_0198_),
    .A2(_1248_),
    .B(_1270_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2495_ (.A1(_0202_),
    .A2(_1297_),
    .B(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2496_ (.I(_0207_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2497_ (.A1(_1264_),
    .A2(_0239_),
    .A3(_1274_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2498_ (.A1(_0198_),
    .A2(_1274_),
    .B(_0202_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2499_ (.A1(_0245_),
    .A2(_1362_),
    .B(_0246_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(_0244_),
    .A2(_0247_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2501_ (.A1(_1256_),
    .A2(_0243_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2502_ (.A1(_0243_),
    .A2(_0249_),
    .B(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2503_ (.A1(_1341_),
    .A2(_0241_),
    .B1(_0251_),
    .B2(_0122_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2504_ (.I0(_0549_),
    .I1(_0189_),
    .S(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2505_ (.A1(_0238_),
    .A2(_0253_),
    .B(_0128_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2506_ (.A1(_0073_),
    .A2(_0086_),
    .A3(_0146_),
    .A4(_0210_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_0552_),
    .A2(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2508_ (.I(_1324_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2509_ (.A1(_1336_),
    .A2(_0058_),
    .B1(_0182_),
    .B2(_0174_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2510_ (.A1(_0180_),
    .A2(_1289_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2511_ (.A1(_1301_),
    .A2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2512_ (.A1(_0182_),
    .A2(_0261_),
    .B(_1276_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2513_ (.A1(_0257_),
    .A2(_0258_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2514_ (.A1(_0256_),
    .A2(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2515_ (.I(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2516_ (.I(_0144_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2517_ (.A1(_1243_),
    .A2(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2518_ (.A1(_1250_),
    .A2(_1289_),
    .B1(_0159_),
    .B2(_1340_),
    .C(_1242_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2519_ (.A1(_1324_),
    .A2(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2520_ (.A1(_1230_),
    .A2(_1297_),
    .B(_0054_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2521_ (.A1(_0098_),
    .A2(_0271_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2522_ (.A1(_0267_),
    .A2(_0269_),
    .B(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2523_ (.A1(_0213_),
    .A2(_0220_),
    .B(_0026_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2524_ (.A1(_0273_),
    .A2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2525_ (.A1(_0041_),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2526_ (.A1(_0254_),
    .A2(_0265_),
    .A3(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2527_ (.A1(_0236_),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2528_ (.A1(_0236_),
    .A2(_0277_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2529_ (.A1(_0278_),
    .A2(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2530_ (.A1(_0224_),
    .A2(_0229_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2531_ (.A1(_0230_),
    .A2(_0233_),
    .B(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2532_ (.A1(_0280_),
    .A2(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2533_ (.I(_0284_),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2534_ (.A1(_0114_),
    .A2(_0126_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2535_ (.A1(_0285_),
    .A2(_0252_),
    .B(net44),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2536_ (.I(_0257_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2537_ (.I(_0244_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2538_ (.A1(_0288_),
    .A2(_0117_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2539_ (.A1(_0239_),
    .A2(_0179_),
    .A3(_0180_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2540_ (.I(_1266_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2541_ (.A1(_0292_),
    .A2(_0302_),
    .B(_1330_),
    .C(_0120_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2542_ (.A1(_0290_),
    .A2(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2543_ (.A1(_0289_),
    .A2(_0266_),
    .B(_0294_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2544_ (.A1(_1348_),
    .A2(_0260_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2545_ (.A1(_0194_),
    .A2(_0141_),
    .B(_0240_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2546_ (.A1(_0141_),
    .A2(_0296_),
    .B(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2547_ (.A1(_0287_),
    .A2(_0295_),
    .B(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2548_ (.A1(_0286_),
    .A2(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2549_ (.A1(_0238_),
    .A2(_0300_),
    .B(_0226_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2550_ (.I(_0026_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2551_ (.A1(_0213_),
    .A2(_0220_),
    .A3(_0273_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2552_ (.A1(_0303_),
    .A2(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2553_ (.I(_1272_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2554_ (.A1(_0207_),
    .A2(_0306_),
    .A3(_1330_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2555_ (.A1(_0120_),
    .A2(_0197_),
    .B(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2556_ (.A1(_0138_),
    .A2(_0078_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2557_ (.A1(_0203_),
    .A2(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2558_ (.I0(_0307_),
    .I1(_0308_),
    .S(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2559_ (.A1(_0054_),
    .A2(_0240_),
    .B1(_0311_),
    .B2(_0257_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2560_ (.A1(_0305_),
    .A2(_0312_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2561_ (.A1(_0041_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2562_ (.A1(_1367_),
    .A2(_0052_),
    .B(_0058_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(_0257_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2564_ (.I(_0202_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2565_ (.A1(_0318_),
    .A2(_0292_),
    .B(_0244_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2566_ (.A1(_0317_),
    .A2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2567_ (.A1(_0149_),
    .A2(_0247_),
    .B1(_0316_),
    .B2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2568_ (.A1(_0255_),
    .A2(_0263_),
    .B(_0552_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2569_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2570_ (.A1(_0546_),
    .A2(_0321_),
    .B(_0323_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2571_ (.A1(_0315_),
    .A2(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2572_ (.A1(_0301_),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2573_ (.A1(_0265_),
    .A2(_0276_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2574_ (.A1(_0265_),
    .A2(_0276_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2575_ (.A1(_0254_),
    .A2(_0328_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2576_ (.A1(_0327_),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2577_ (.A1(_0230_),
    .A2(_0233_),
    .B(_0279_),
    .C(_0282_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2578_ (.A1(_0278_),
    .A2(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2579_ (.A1(_0331_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2580_ (.I(_0334_),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2581_ (.A1(_0315_),
    .A2(_0325_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2582_ (.I(_0326_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2583_ (.A1(_0301_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2584_ (.A1(_0114_),
    .A2(_0071_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2585_ (.A1(_0238_),
    .A2(_0338_),
    .B(_0021_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2586_ (.I(_0130_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2587_ (.I(_0318_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2588_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2589_ (.A1(_0342_),
    .A2(_1303_),
    .B1(_0154_),
    .B2(_0206_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2590_ (.I(_0288_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2591_ (.A1(_0184_),
    .A2(_0266_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2592_ (.I(_0317_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2593_ (.A1(_0345_),
    .A2(_0346_),
    .B(_0067_),
    .C(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2594_ (.I(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2595_ (.A1(_0341_),
    .A2(_0117_),
    .A3(_0154_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2596_ (.A1(_0342_),
    .A2(_0139_),
    .B(_0350_),
    .C(_1371_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2597_ (.A1(_1344_),
    .A2(_0343_),
    .B(_0349_),
    .C(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2598_ (.I(_0286_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2599_ (.A1(_0353_),
    .A2(_0352_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2600_ (.A1(_0549_),
    .A2(_0352_),
    .B(_0354_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2601_ (.A1(_0340_),
    .A2(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2602_ (.A1(_0339_),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2603_ (.A1(_0341_),
    .A2(_0089_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2604_ (.A1(_0287_),
    .A2(_0197_),
    .A3(_0068_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2605_ (.A1(_0194_),
    .A2(_1351_),
    .A3(_1330_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2606_ (.A1(_0359_),
    .A2(_0360_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2607_ (.A1(_0322_),
    .A2(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2608_ (.I(_0317_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2609_ (.I(_0174_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2610_ (.A1(_0365_),
    .A2(_0204_),
    .A3(_0078_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2611_ (.A1(_0055_),
    .A2(_0319_),
    .B1(_0367_),
    .B2(_0206_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2612_ (.A1(_0364_),
    .A2(_0368_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2613_ (.I(_0212_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2614_ (.A1(_0305_),
    .A2(_0369_),
    .B(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2615_ (.A1(_0305_),
    .A2(_0369_),
    .B(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2616_ (.A1(_0363_),
    .A2(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2617_ (.A1(_0358_),
    .A2(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2618_ (.A1(_0335_),
    .A2(_0337_),
    .B(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2619_ (.I(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2620_ (.A1(_0335_),
    .A2(_0337_),
    .A3(_0374_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(_0376_),
    .A2(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2622_ (.A1(_0327_),
    .A2(_0330_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2623_ (.A1(_0278_),
    .A2(_0332_),
    .A3(_0331_),
    .B(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2624_ (.A1(_0379_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2625_ (.I(_0382_),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2626_ (.I(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2627_ (.A1(_1371_),
    .A2(_0203_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2628_ (.A1(_0318_),
    .A2(_0288_),
    .A3(_1346_),
    .A4(_0154_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2629_ (.A1(_1334_),
    .A2(_0198_),
    .B(_0179_),
    .C(_0203_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2630_ (.A1(_0059_),
    .A2(_0386_),
    .B(_0365_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2631_ (.A1(_0287_),
    .A2(_0385_),
    .A3(_0388_),
    .B1(_0116_),
    .B2(_0350_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2632_ (.A1(_0242_),
    .A2(_0384_),
    .B(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2633_ (.I0(_0383_),
    .I1(_0353_),
    .S(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2634_ (.A1(_0340_),
    .A2(_0391_),
    .B(_0192_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2635_ (.A1(_0184_),
    .A2(_0266_),
    .B1(_0176_),
    .B2(_0309_),
    .C(_0244_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2636_ (.A1(_0255_),
    .A2(_0263_),
    .A3(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2637_ (.A1(_1367_),
    .A2(_1371_),
    .B(_1283_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2638_ (.A1(_0395_),
    .A2(_0546_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2639_ (.A1(_0248_),
    .A2(\p_shaping_I.p_shaping_I.bit_in ),
    .A3(_0394_),
    .B1(_0396_),
    .B2(_0107_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2640_ (.I(_0303_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2641_ (.A1(_0174_),
    .A2(_1310_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2642_ (.A1(_0400_),
    .A2(_0206_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2643_ (.I(_0182_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2644_ (.A1(_0292_),
    .A2(_1235_),
    .B(_0318_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2645_ (.A1(_0075_),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2646_ (.A1(_0402_),
    .A2(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2647_ (.A1(_0365_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2648_ (.A1(_0401_),
    .A2(_0406_),
    .B(_0317_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2649_ (.A1(_0178_),
    .A2(_0213_),
    .A3(_0220_),
    .A4(_0273_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2650_ (.A1(_0303_),
    .A2(_0408_),
    .B(_0407_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2651_ (.A1(_0399_),
    .A2(_0407_),
    .B(_0410_),
    .C(_0370_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2652_ (.A1(_0397_),
    .A2(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2653_ (.A1(_0392_),
    .A2(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2654_ (.A1(_0339_),
    .A2(_0357_),
    .A3(_0373_),
    .B1(_0372_),
    .B2(_0363_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2655_ (.A1(_0413_),
    .A2(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2656_ (.A1(_0375_),
    .A2(_0381_),
    .B(_0378_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2657_ (.A1(_0415_),
    .A2(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2658_ (.I(_0417_),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2659_ (.A1(_0397_),
    .A2(_0411_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2660_ (.A1(_0392_),
    .A2(_0412_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2661_ (.A1(_0288_),
    .A2(_0117_),
    .A3(_0403_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2662_ (.A1(_0197_),
    .A2(_0421_),
    .B(_0400_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2663_ (.A1(_0287_),
    .A2(_0393_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2664_ (.A1(_0364_),
    .A2(_0422_),
    .B(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2665_ (.I0(_0353_),
    .I1(_0383_),
    .S(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2666_ (.A1(_0340_),
    .A2(_0425_),
    .B(_0192_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2667_ (.A1(_0255_),
    .A2(_0263_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2668_ (.A1(\p_shaping_I.p_shaping_I.bit_in ),
    .A2(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2669_ (.A1(_0364_),
    .A2(_1328_),
    .A3(_0054_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2670_ (.A1(_0395_),
    .A2(_0429_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2671_ (.I0(\p_shaping_I.p_shaping_I.bit_in ),
    .I1(_0428_),
    .S(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2672_ (.A1(_0341_),
    .A2(_0306_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2673_ (.A1(_0179_),
    .A2(_1347_),
    .A3(_0306_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2674_ (.A1(_0345_),
    .A2(_0433_),
    .B1(_0319_),
    .B2(_0434_),
    .C(_0364_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2675_ (.I0(_0305_),
    .I1(_0399_),
    .S(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2676_ (.A1(_0370_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2677_ (.A1(_0426_),
    .A2(_0432_),
    .A3(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2678_ (.A1(_0418_),
    .A2(_0420_),
    .B(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2679_ (.A1(_0418_),
    .A2(_0420_),
    .A3(_0438_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2680_ (.A1(_0439_),
    .A2(_0440_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2681_ (.A1(_0413_),
    .A2(_0414_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2682_ (.A1(_0415_),
    .A2(_0416_),
    .B(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2683_ (.A1(_0442_),
    .A2(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2684_ (.I(_0445_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2685_ (.A1(_0415_),
    .A2(_0442_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2686_ (.A1(_0375_),
    .A2(_0381_),
    .B(_0446_),
    .C(_0378_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2687_ (.A1(_0443_),
    .A2(_0439_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2688_ (.A1(_0440_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2689_ (.A1(_0395_),
    .A2(_0322_),
    .B(_0396_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2690_ (.A1(_0306_),
    .A2(_1316_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2691_ (.A1(_0345_),
    .A2(_0433_),
    .B(_0452_),
    .C(_0347_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2692_ (.A1(_0399_),
    .A2(_0304_),
    .B(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2693_ (.A1(_0399_),
    .A2(_0453_),
    .B(_0454_),
    .C(_0370_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2694_ (.A1(_0450_),
    .A2(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2695_ (.A1(_0342_),
    .A2(_1297_),
    .B(_0319_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2696_ (.A1(_1344_),
    .A2(_0271_),
    .B1(_0457_),
    .B2(_0347_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2697_ (.A1(_0050_),
    .A2(_0338_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2698_ (.A1(_0238_),
    .A2(_0353_),
    .B(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2699_ (.A1(_0458_),
    .A2(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2700_ (.A1(_1279_),
    .A2(_0461_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2701_ (.A1(_0456_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2702_ (.A1(_0432_),
    .A2(_0437_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2703_ (.A1(_0426_),
    .A2(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2704_ (.A1(_0432_),
    .A2(_0437_),
    .B(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2705_ (.A1(_0464_),
    .A2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2706_ (.A1(_0447_),
    .A2(_0449_),
    .B(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2707_ (.A1(_0468_),
    .A2(_0447_),
    .A3(_0449_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2708_ (.A1(_0469_),
    .A2(_0470_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2709_ (.A1(_0450_),
    .A2(_0455_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2710_ (.A1(_0456_),
    .A2(_0463_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2711_ (.I(_0342_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2712_ (.A1(_0474_),
    .A2(_0240_),
    .B(_1299_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2713_ (.A1(_0285_),
    .A2(_0252_),
    .B(_0475_),
    .C(_0383_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2714_ (.A1(_0383_),
    .A2(_0475_),
    .B(_0476_),
    .C(_0340_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2715_ (.A1(_0226_),
    .A2(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2716_ (.A1(_0456_),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2717_ (.A1(_0471_),
    .A2(_0473_),
    .B(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2718_ (.A1(_0471_),
    .A2(_0473_),
    .A3(_0479_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2719_ (.A1(_0480_),
    .A2(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(_0464_),
    .A2(_0467_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2721_ (.A1(_0484_),
    .A2(_0469_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2722_ (.A1(_0482_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2723_ (.I(_0486_),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2724_ (.A1(_0484_),
    .A2(_0469_),
    .A3(_0480_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2725_ (.A1(_1279_),
    .A2(_0460_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2726_ (.A1(_0450_),
    .A2(_0455_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2727_ (.A1(_0489_),
    .A2(_0478_),
    .B(_0471_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2728_ (.A1(_0488_),
    .A2(_0490_),
    .B(_0481_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2729_ (.A1(_0488_),
    .A2(_0490_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2730_ (.A1(_0487_),
    .A2(_0491_),
    .B(_0492_),
    .ZN(net9));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2731_ (.A1(_0040_),
    .A2(_0044_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2732_ (.I(_0494_),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2733_ (.A1(\p_shaping_Q.p_shaping_I.counter[0] ),
    .A2(_0756_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2734_ (.A1(_0007_),
    .A2(_0495_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2735_ (.A1(net69),
    .A2(net3),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2736_ (.I(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2737_ (.A1(_0239_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2738_ (.I(_0498_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2739_ (.I(_0496_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2740_ (.I(_0499_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2741_ (.A1(_0550_),
    .A2(_1226_),
    .B(_0497_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2742_ (.A1(_1334_),
    .A2(_0501_),
    .B(_0502_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2743_ (.A1(_0292_),
    .A2(_0501_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2744_ (.A1(_0089_),
    .A2(_0501_),
    .B(_0503_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2745_ (.A1(_1347_),
    .A2(_0496_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2746_ (.A1(_0474_),
    .A2(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2747_ (.I(_0505_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2748_ (.A1(_0550_),
    .A2(_0497_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2749_ (.A1(_0474_),
    .A2(_0345_),
    .A3(_0504_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2750_ (.A1(_0474_),
    .A2(_0504_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2751_ (.A1(_0365_),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2752_ (.A1(_0507_),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2753_ (.A1(_0506_),
    .A2(_0511_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2754_ (.A1(_0347_),
    .A2(_0507_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2755_ (.A1(_0506_),
    .A2(_0512_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2756_ (.A1(_0906_),
    .A2(_0499_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2757_ (.I(_0513_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2758_ (.A1(_0591_),
    .A2(_0497_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2759_ (.A1(net50),
    .A2(_1007_),
    .A3(_0501_),
    .B(_0514_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2760_ (.A1(_0913_),
    .A2(_0499_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2761_ (.A1(_1045_),
    .A2(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2762_ (.I(_0517_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2763_ (.A1(_0818_),
    .A2(_0913_),
    .A3(_0496_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2764_ (.A1(_1145_),
    .A2(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2765_ (.I(_0519_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2766_ (.A1(_1145_),
    .A2(_1051_),
    .A3(_0518_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2767_ (.A1(_1145_),
    .A2(_0518_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2768_ (.A1(_0870_),
    .A2(_0540_),
    .A3(_0499_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2769_ (.A1(_1119_),
    .A2(_0521_),
    .B(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2770_ (.A1(_0520_),
    .A2(_0523_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2771_ (.I(_0525_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2772_ (.A1(_1117_),
    .A2(_0520_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2773_ (.A1(_0522_),
    .A2(_0526_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2774_ (.A1(_0041_),
    .A2(\p_shaping_I.p_shaping_I.counter[0] ),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2775_ (.A1(_0021_),
    .A2(_0527_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2776_ (.D(_0006_),
    .RN(net61),
    .CLK(net48),
    .Q(\p_shaping_Q.p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2777_ (.D(_0007_),
    .RN(net61),
    .CLK(net49),
    .Q(\p_shaping_Q.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2778_ (.D(\gen_sym.Reg_2M.data_in ),
    .RN(net59),
    .CLK(net45),
    .Q(\gen_sym.Reg_Sym.data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2779_ (.D(\gen_sym.Reg_2M.data_out ),
    .RN(net60),
    .CLK(net45),
    .Q(\gen_sym.Reg_Sym.data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2780_ (.D(\gen_sym.Reg_2M.data_in ),
    .RN(net59),
    .CLK(\gen_sym.Reg_2M.enable ),
    .Q(\gen_sym.Reg_2M.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2781_ (.D(\mapper.bit_Q[1] ),
    .RN(net60),
    .CLK(net49),
    .Q(\p_shaping_Q.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2782_ (.D(net44),
    .RN(net64),
    .CLK(net45),
    .Q(\p_shaping_I.p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2783_ (.D(_0000_),
    .Q(\p_shaping_I.p_shaping_I.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2784_ (.D(_0008_),
    .RN(net57),
    .CLK(net68),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2785_ (.D(_0009_),
    .RN(net56),
    .CLK(net66),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2786_ (.D(_0010_),
    .RN(net56),
    .CLK(net67),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2787_ (.D(_0011_),
    .RN(net58),
    .CLK(net69),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _2788_ (.D(_0012_),
    .RN(net59),
    .CLK(net70),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2789_ (.D(_0013_),
    .RN(net59),
    .CLK(net70),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2790_ (.D(\p_shaping_I.p_shaping_I.bit_in ),
    .RN(net63),
    .CLK(net46),
    .Q(\p_shaping_I.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2791_ (.D(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .RN(net61),
    .CLK(net48),
    .Q(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2792_ (.D(_0002_),
    .Q(\p_shaping_Q.p_shaping_I.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 _2793_ (.D(_0014_),
    .SETN(net55),
    .CLK(net66),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2794_ (.D(_0015_),
    .RN(net55),
    .CLK(net67),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2795_ (.D(_0016_),
    .RN(net55),
    .CLK(net66),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 _2796_ (.D(_0017_),
    .SETN(net55),
    .CLK(net66),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 _2797_ (.D(_0018_),
    .SETN(net57),
    .CLK(net68),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2798_ (.D(_0019_),
    .RN(net58),
    .CLK(net69),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2799_ (.D(\p_shaping_Q.p_shaping_I.bit_in ),
    .RN(net60),
    .CLK(net49),
    .Q(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2800_ (.D(_0020_),
    .RN(net62),
    .CLK(net47),
    .Q(\p_shaping_I.p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2801_ (.D(_0021_),
    .RN(net62),
    .CLK(net47),
    .Q(\p_shaping_I.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout44 (.I(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout46 (.I(_0004_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout47 (.I(_0004_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout50 (.I(_0005_),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout51 (.I(net43),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout52 (.I(net40),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout53 (.I(net37),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout54 (.I(net34),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout55 (.I(net57),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout58 (.I(net65),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout59 (.I(net64),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout60 (.I(net63),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout61 (.I(net63),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout62 (.I(net63),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout63 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout65 (.I(net5),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout66 (.I(net68),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout68 (.I(net69),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout69 (.I(net4),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout70 (.I(net4),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(ACK),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(Bit_In),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(EN),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(REQ_SAMPLE),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(RST),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output10 (.I(net10),
    .Z(I[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output11 (.I(net11),
    .Z(I[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output12 (.I(net12),
    .Z(I[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(I[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(I[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net15),
    .Z(I[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(I[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(I[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(I[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(Q[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(Q[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(Q[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(Q[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(Q[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(Q[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(Q[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(Q[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(Q[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(Q[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(Q[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output30 (.I(net30),
    .Z(Q[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output31 (.I(net31),
    .Z(Q[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output32 (.I(net32),
    .Z(addI[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output33 (.I(net33),
    .Z(addI[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output34 (.I(net54),
    .Z(addI[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output35 (.I(net35),
    .Z(addI[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output36 (.I(net36),
    .Z(addI[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output37 (.I(net37),
    .Z(addI[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output38 (.I(net38),
    .Z(addQ[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output39 (.I(net39),
    .Z(addQ[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output40 (.I(net52),
    .Z(addQ[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output41 (.I(net41),
    .Z(addQ[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output42 (.I(net42),
    .Z(addQ[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output43 (.I(net51),
    .Z(addQ[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(I[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(I[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(I[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output9 (.I(net9),
    .Z(I[12]));
 assign io_oeb[0] = net100;
 assign io_oeb[10] = net72;
 assign io_oeb[11] = net73;
 assign io_oeb[12] = net74;
 assign io_oeb[13] = net75;
 assign io_oeb[14] = net76;
 assign io_oeb[15] = net77;
 assign io_oeb[16] = net78;
 assign io_oeb[17] = net79;
 assign io_oeb[18] = net80;
 assign io_oeb[19] = net81;
 assign io_oeb[1] = net101;
 assign io_oeb[20] = net82;
 assign io_oeb[21] = net83;
 assign io_oeb[22] = net84;
 assign io_oeb[23] = net85;
 assign io_oeb[24] = net86;
 assign io_oeb[25] = net87;
 assign io_oeb[26] = net88;
 assign io_oeb[27] = net89;
 assign io_oeb[28] = net90;
 assign io_oeb[29] = net91;
 assign io_oeb[2] = net102;
 assign io_oeb[30] = net92;
 assign io_oeb[31] = net93;
 assign io_oeb[32] = net94;
 assign io_oeb[33] = net95;
 assign io_oeb[34] = net96;
 assign io_oeb[35] = net97;
 assign io_oeb[36] = net98;
 assign io_oeb[37] = net99;
 assign io_oeb[3] = net103;
 assign io_oeb[4] = net104;
 assign io_oeb[5] = net105;
 assign io_oeb[6] = net106;
 assign io_oeb[7] = net107;
 assign io_oeb[8] = net108;
 assign io_oeb[9] = net71;
endmodule

